


module picorv32_pads(clk, resetn, trap, mem_valid, mem_instr, mem_ready,
     mem_addr, mem_wdata, mem_wstrb, mem_rdata, mem_la_read,
     mem_la_write, mem_la_addr, mem_la_wdata, mem_la_wstrb, pcpi_valid,
     pcpi_insn, pcpi_rs1, pcpi_rs2, pcpi_wr, pcpi_rd, pcpi_wait,
     pcpi_ready, irq, eoi, trace_valid, trace_data, 
     clk_w, resetn_w, trap_w, mem_valid_w, mem_instr_w, mem_ready_w,
     mem_addr_w, mem_wdata_w, mem_wstrb_w, mem_rdata_w, mem_la_read_w,
     mem_la_write_w, mem_la_addr_w, mem_la_wdata_w, mem_la_wstrb_w, pcpi_valid_w,
     pcpi_insn_w, pcpi_rs1_w, pcpi_rs2_w, pcpi_wr_w, pcpi_rd_w, pcpi_wait_w,
     pcpi_ready_w, irq_w, eoi_w, trace_valid_w, trace_data_w, VSS, VDD);

     input clk, resetn, mem_ready, pcpi_wr, pcpi_wait, pcpi_ready;
     input [31:0] mem_rdata, pcpi_rd, irq;
     output trap, mem_valid, mem_instr, mem_la_read, mem_la_write,
          pcpi_valid, trace_valid;
     output [31:0] mem_addr, mem_wdata, mem_la_addr, mem_la_wdata,
          pcpi_insn, pcpi_rs1, pcpi_rs2, eoi;
     output [3:0] mem_wstrb, mem_la_wstrb;
     output [35:0] trace_data;

     output clk_w, resetn_w, mem_ready_w, pcpi_wr_w, pcpi_wait_w, pcpi_ready_w;
     output [31:0] mem_rdata_w, pcpi_rd_w, irq_w;
     input trap_w, mem_valid_w, mem_instr_w, mem_la_read_w, mem_la_write_w,
          pcpi_valid_w, trace_valid_w;
     input [31:0] mem_addr_w, mem_wdata_w, mem_la_addr_w, mem_la_wdata_w,
          pcpi_insn_w, pcpi_rs1_w, pcpi_rs2_w, eoi_w;
     input [3:0] mem_wstrb_w, mem_la_wstrb_w;
     input [35:0] trace_data_w;

     wire clk, resetn, mem_ready, pcpi_wr, pcpi_wait, pcpi_ready;
     wire [31:0] mem_rdata, pcpi_rd, irq;
     wire trap, mem_valid, mem_instr, mem_la_read, mem_la_write,
          pcpi_valid, trace_valid;
     wire [31:0] mem_addr, mem_wdata, mem_la_addr, mem_la_wdata,
          pcpi_insn, pcpi_rs1, pcpi_rs2, eoi;
     wire [3:0] mem_wstrb, mem_la_wstrb;
     wire [35:0] trace_data;


     input VSS, VDD;
     supply0 VSS;
     supply1 VDD;

     
//Insert Pads
PADVSS pad_vss(.VSS(VSS), .VDD(VDD), .VDDIOR(VDD), .VSSIOR(VSS));  
PADVDD pad_vdd(.VSS(VSS), .VDD(VDD), .VDDIOR(VDD), .VSSIOR(VSS));
PADDI pad_clk(.PAD(clk), .Y(clk_w), .VDD(VDD), .VSS(VSS));
PADDI pad_resetn(.PAD(resetn), .Y(resetn_w), .VDD(VDD), .VSS(VSS));
PADDI pad_mem_ready(.PAD(mem_ready), .Y(mem_ready_w), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_wr(.PAD(pcpi_wr), .Y(pcpi_wr_w), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_wait(.PAD(pcpi_wait), .Y(pcpi_wait_w), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_ready(.PAD(pcpi_ready), .Y(pcpi_ready_w), .VDD(VDD), .VSS(VSS));
PADDO pad_trap(.PAD(trap), .A(trap_w), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_valid(.PAD(mem_valid), .A(mem_valid_w), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_instr(.PAD(mem_instr), .A(mem_instr_w), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_read(.PAD(mem_la_read), .A(mem_la_read_w), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_write(.PAD(mem_la_write), .A(mem_la_write_w), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_valid(.PAD(pcpi_valid), .A(pcpi_valid_w), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_valid(.PAD(trace_valid), .A(trace_valid_w), .VDD(VDD), .VSS(VSS));
PADDI pad_mem_rdata0(.PAD(mem_rdata[0]), .Y(mem_rdata_w[0]), .VDD(VDD), .VSS(VSS));
PADDI pad_mem_rdata1(.PAD(mem_rdata[1]), .Y(mem_rdata_w[1]), .VDD(VDD), .VSS(VSS));
PADDI pad_mem_rdata2(.PAD(mem_rdata[2]), .Y(mem_rdata_w[2]), .VDD(VDD), .VSS(VSS));
PADDI pad_mem_rdata3(.PAD(mem_rdata[3]), .Y(mem_rdata_w[3]), .VDD(VDD), .VSS(VSS));
PADDI pad_mem_rdata4(.PAD(mem_rdata[4]), .Y(mem_rdata_w[4]), .VDD(VDD), .VSS(VSS));
PADDI pad_mem_rdata5(.PAD(mem_rdata[5]), .Y(mem_rdata_w[5]), .VDD(VDD), .VSS(VSS));
PADDI pad_mem_rdata6(.PAD(mem_rdata[6]), .Y(mem_rdata_w[6]), .VDD(VDD), .VSS(VSS));
PADDI pad_mem_rdata7(.PAD(mem_rdata[7]), .Y(mem_rdata_w[7]), .VDD(VDD), .VSS(VSS));
PADDI pad_mem_rdata8(.PAD(mem_rdata[8]), .Y(mem_rdata_w[8]), .VDD(VDD), .VSS(VSS));
PADDI pad_mem_rdata9(.PAD(mem_rdata[9]), .Y(mem_rdata_w[9]), .VDD(VDD), .VSS(VSS));
PADDI pad_mem_rdata10(.PAD(mem_rdata[10]), .Y(mem_rdata_w[10]), .VDD(VDD), .VSS(VSS));
PADDI pad_mem_rdata11(.PAD(mem_rdata[11]), .Y(mem_rdata_w[11]), .VDD(VDD), .VSS(VSS));
PADDI pad_mem_rdata12(.PAD(mem_rdata[12]), .Y(mem_rdata_w[12]), .VDD(VDD), .VSS(VSS));
PADDI pad_mem_rdata13(.PAD(mem_rdata[13]), .Y(mem_rdata_w[13]), .VDD(VDD), .VSS(VSS));
PADDI pad_mem_rdata14(.PAD(mem_rdata[14]), .Y(mem_rdata_w[14]), .VDD(VDD), .VSS(VSS));
PADDI pad_mem_rdata15(.PAD(mem_rdata[15]), .Y(mem_rdata_w[15]), .VDD(VDD), .VSS(VSS));
PADDI pad_mem_rdata16(.PAD(mem_rdata[16]), .Y(mem_rdata_w[16]), .VDD(VDD), .VSS(VSS));
PADDI pad_mem_rdata17(.PAD(mem_rdata[17]), .Y(mem_rdata_w[17]), .VDD(VDD), .VSS(VSS));
PADDI pad_mem_rdata18(.PAD(mem_rdata[18]), .Y(mem_rdata_w[18]), .VDD(VDD), .VSS(VSS));
PADDI pad_mem_rdata19(.PAD(mem_rdata[19]), .Y(mem_rdata_w[19]), .VDD(VDD), .VSS(VSS));
PADDI pad_mem_rdata20(.PAD(mem_rdata[20]), .Y(mem_rdata_w[20]), .VDD(VDD), .VSS(VSS));
PADDI pad_mem_rdata21(.PAD(mem_rdata[21]), .Y(mem_rdata_w[21]), .VDD(VDD), .VSS(VSS));
PADDI pad_mem_rdata22(.PAD(mem_rdata[22]), .Y(mem_rdata_w[22]), .VDD(VDD), .VSS(VSS));
PADDI pad_mem_rdata23(.PAD(mem_rdata[23]), .Y(mem_rdata_w[23]), .VDD(VDD), .VSS(VSS));
PADDI pad_mem_rdata24(.PAD(mem_rdata[24]), .Y(mem_rdata_w[24]), .VDD(VDD), .VSS(VSS));
PADDI pad_mem_rdata25(.PAD(mem_rdata[25]), .Y(mem_rdata_w[25]), .VDD(VDD), .VSS(VSS));
PADDI pad_mem_rdata26(.PAD(mem_rdata[26]), .Y(mem_rdata_w[26]), .VDD(VDD), .VSS(VSS));
PADDI pad_mem_rdata27(.PAD(mem_rdata[27]), .Y(mem_rdata_w[27]), .VDD(VDD), .VSS(VSS));
PADDI pad_mem_rdata28(.PAD(mem_rdata[28]), .Y(mem_rdata_w[28]), .VDD(VDD), .VSS(VSS));
PADDI pad_mem_rdata29(.PAD(mem_rdata[29]), .Y(mem_rdata_w[29]), .VDD(VDD), .VSS(VSS));
PADDI pad_mem_rdata30(.PAD(mem_rdata[30]), .Y(mem_rdata_w[30]), .VDD(VDD), .VSS(VSS));
PADDI pad_mem_rdata31(.PAD(mem_rdata[31]), .Y(mem_rdata_w[31]), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_rd0(.PAD(pcpi_rd[0]), .Y(pcpi_rd_w[0]), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_rd1(.PAD(pcpi_rd[1]), .Y(pcpi_rd_w[1]), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_rd2(.PAD(pcpi_rd[2]), .Y(pcpi_rd_w[2]), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_rd3(.PAD(pcpi_rd[3]), .Y(pcpi_rd_w[3]), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_rd4(.PAD(pcpi_rd[4]), .Y(pcpi_rd_w[4]), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_rd5(.PAD(pcpi_rd[5]), .Y(pcpi_rd_w[5]), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_rd6(.PAD(pcpi_rd[6]), .Y(pcpi_rd_w[6]), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_rd7(.PAD(pcpi_rd[7]), .Y(pcpi_rd_w[7]), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_rd8(.PAD(pcpi_rd[8]), .Y(pcpi_rd_w[8]), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_rd9(.PAD(pcpi_rd[9]), .Y(pcpi_rd_w[9]), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_rd10(.PAD(pcpi_rd[10]), .Y(pcpi_rd_w[10]), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_rd11(.PAD(pcpi_rd[11]), .Y(pcpi_rd_w[11]), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_rd12(.PAD(pcpi_rd[12]), .Y(pcpi_rd_w[12]), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_rd13(.PAD(pcpi_rd[13]), .Y(pcpi_rd_w[13]), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_rd14(.PAD(pcpi_rd[14]), .Y(pcpi_rd_w[14]), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_rd15(.PAD(pcpi_rd[15]), .Y(pcpi_rd_w[15]), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_rd16(.PAD(pcpi_rd[16]), .Y(pcpi_rd_w[16]), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_rd17(.PAD(pcpi_rd[17]), .Y(pcpi_rd_w[17]), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_rd18(.PAD(pcpi_rd[18]), .Y(pcpi_rd_w[18]), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_rd19(.PAD(pcpi_rd[19]), .Y(pcpi_rd_w[19]), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_rd20(.PAD(pcpi_rd[20]), .Y(pcpi_rd_w[20]), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_rd21(.PAD(pcpi_rd[21]), .Y(pcpi_rd_w[21]), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_rd22(.PAD(pcpi_rd[22]), .Y(pcpi_rd_w[22]), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_rd23(.PAD(pcpi_rd[23]), .Y(pcpi_rd_w[23]), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_rd24(.PAD(pcpi_rd[24]), .Y(pcpi_rd_w[24]), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_rd25(.PAD(pcpi_rd[25]), .Y(pcpi_rd_w[25]), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_rd26(.PAD(pcpi_rd[26]), .Y(pcpi_rd_w[26]), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_rd27(.PAD(pcpi_rd[27]), .Y(pcpi_rd_w[27]), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_rd28(.PAD(pcpi_rd[28]), .Y(pcpi_rd_w[28]), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_rd29(.PAD(pcpi_rd[29]), .Y(pcpi_rd_w[29]), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_rd30(.PAD(pcpi_rd[30]), .Y(pcpi_rd_w[30]), .VDD(VDD), .VSS(VSS));
PADDI pad_pcpi_rd31(.PAD(pcpi_rd[31]), .Y(pcpi_rd_w[31]), .VDD(VDD), .VSS(VSS));
PADDI pad_irq0(.PAD(irq[0]), .Y(irq_w[0]), .VDD(VDD), .VSS(VSS));
PADDI pad_irq1(.PAD(irq[1]), .Y(irq_w[1]), .VDD(VDD), .VSS(VSS));
PADDI pad_irq2(.PAD(irq[2]), .Y(irq_w[2]), .VDD(VDD), .VSS(VSS));
PADDI pad_irq3(.PAD(irq[3]), .Y(irq_w[3]), .VDD(VDD), .VSS(VSS));
PADDI pad_irq4(.PAD(irq[4]), .Y(irq_w[4]), .VDD(VDD), .VSS(VSS));
PADDI pad_irq5(.PAD(irq[5]), .Y(irq_w[5]), .VDD(VDD), .VSS(VSS));
PADDI pad_irq6(.PAD(irq[6]), .Y(irq_w[6]), .VDD(VDD), .VSS(VSS));
PADDI pad_irq7(.PAD(irq[7]), .Y(irq_w[7]), .VDD(VDD), .VSS(VSS));
PADDI pad_irq8(.PAD(irq[8]), .Y(irq_w[8]), .VDD(VDD), .VSS(VSS));
PADDI pad_irq9(.PAD(irq[9]), .Y(irq_w[9]), .VDD(VDD), .VSS(VSS));
PADDI pad_irq10(.PAD(irq[10]), .Y(irq_w[10]), .VDD(VDD), .VSS(VSS));
PADDI pad_irq11(.PAD(irq[11]), .Y(irq_w[11]), .VDD(VDD), .VSS(VSS));
PADDI pad_irq12(.PAD(irq[12]), .Y(irq_w[12]), .VDD(VDD), .VSS(VSS));
PADDI pad_irq13(.PAD(irq[13]), .Y(irq_w[13]), .VDD(VDD), .VSS(VSS));
PADDI pad_irq14(.PAD(irq[14]), .Y(irq_w[14]), .VDD(VDD), .VSS(VSS));
PADDI pad_irq15(.PAD(irq[15]), .Y(irq_w[15]), .VDD(VDD), .VSS(VSS));
PADDI pad_irq16(.PAD(irq[16]), .Y(irq_w[16]), .VDD(VDD), .VSS(VSS));
PADDI pad_irq17(.PAD(irq[17]), .Y(irq_w[17]), .VDD(VDD), .VSS(VSS));
PADDI pad_irq18(.PAD(irq[18]), .Y(irq_w[18]), .VDD(VDD), .VSS(VSS));
PADDI pad_irq19(.PAD(irq[19]), .Y(irq_w[19]), .VDD(VDD), .VSS(VSS));
PADDI pad_irq20(.PAD(irq[20]), .Y(irq_w[20]), .VDD(VDD), .VSS(VSS));
PADDI pad_irq21(.PAD(irq[21]), .Y(irq_w[21]), .VDD(VDD), .VSS(VSS));
PADDI pad_irq22(.PAD(irq[22]), .Y(irq_w[22]), .VDD(VDD), .VSS(VSS));
PADDI pad_irq23(.PAD(irq[23]), .Y(irq_w[23]), .VDD(VDD), .VSS(VSS));
PADDI pad_irq24(.PAD(irq[24]), .Y(irq_w[24]), .VDD(VDD), .VSS(VSS));
PADDI pad_irq25(.PAD(irq[25]), .Y(irq_w[25]), .VDD(VDD), .VSS(VSS));
PADDI pad_irq26(.PAD(irq[26]), .Y(irq_w[26]), .VDD(VDD), .VSS(VSS));
PADDI pad_irq27(.PAD(irq[27]), .Y(irq_w[27]), .VDD(VDD), .VSS(VSS));
PADDI pad_irq28(.PAD(irq[28]), .Y(irq_w[28]), .VDD(VDD), .VSS(VSS));
PADDI pad_irq29(.PAD(irq[29]), .Y(irq_w[29]), .VDD(VDD), .VSS(VSS));
PADDI pad_irq30(.PAD(irq[30]), .Y(irq_w[30]), .VDD(VDD), .VSS(VSS));
PADDI pad_irq31(.PAD(irq[31]), .Y(irq_w[31]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_addr0(.PAD(mem_addr[0]), .A(mem_addr_w[0]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_addr1(.PAD(mem_addr[1]), .A(mem_addr_w[1]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_addr2(.PAD(mem_addr[2]), .A(mem_addr_w[2]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_addr3(.PAD(mem_addr[3]), .A(mem_addr_w[3]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_addr4(.PAD(mem_addr[4]), .A(mem_addr_w[4]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_addr5(.PAD(mem_addr[5]), .A(mem_addr_w[5]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_addr6(.PAD(mem_addr[6]), .A(mem_addr_w[6]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_addr7(.PAD(mem_addr[7]), .A(mem_addr_w[7]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_addr8(.PAD(mem_addr[8]), .A(mem_addr_w[8]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_addr9(.PAD(mem_addr[9]), .A(mem_addr_w[9]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_addr10(.PAD(mem_addr[10]), .A(mem_addr_w[10]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_addr11(.PAD(mem_addr[11]), .A(mem_addr_w[11]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_addr12(.PAD(mem_addr[12]), .A(mem_addr_w[12]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_addr13(.PAD(mem_addr[13]), .A(mem_addr_w[13]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_addr14(.PAD(mem_addr[14]), .A(mem_addr_w[14]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_addr15(.PAD(mem_addr[15]), .A(mem_addr_w[15]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_addr16(.PAD(mem_addr[16]), .A(mem_addr_w[16]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_addr17(.PAD(mem_addr[17]), .A(mem_addr_w[17]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_addr18(.PAD(mem_addr[18]), .A(mem_addr_w[18]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_addr19(.PAD(mem_addr[19]), .A(mem_addr_w[19]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_addr20(.PAD(mem_addr[20]), .A(mem_addr_w[20]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_addr21(.PAD(mem_addr[21]), .A(mem_addr_w[21]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_addr22(.PAD(mem_addr[22]), .A(mem_addr_w[22]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_addr23(.PAD(mem_addr[23]), .A(mem_addr_w[23]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_addr24(.PAD(mem_addr[24]), .A(mem_addr_w[24]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_addr25(.PAD(mem_addr[25]), .A(mem_addr_w[25]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_addr26(.PAD(mem_addr[26]), .A(mem_addr_w[26]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_addr27(.PAD(mem_addr[27]), .A(mem_addr_w[27]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_addr28(.PAD(mem_addr[28]), .A(mem_addr_w[28]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_addr29(.PAD(mem_addr[29]), .A(mem_addr_w[29]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_addr30(.PAD(mem_addr[30]), .A(mem_addr_w[30]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_addr31(.PAD(mem_addr[31]), .A(mem_addr_w[31]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wdata0(.PAD(mem_wdata[0]), .A(mem_wdata_w[0]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wdata1(.PAD(mem_wdata[1]), .A(mem_wdata_w[1]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wdata2(.PAD(mem_wdata[2]), .A(mem_wdata_w[2]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wdata3(.PAD(mem_wdata[3]), .A(mem_wdata_w[3]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wdata4(.PAD(mem_wdata[4]), .A(mem_wdata_w[4]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wdata5(.PAD(mem_wdata[5]), .A(mem_wdata_w[5]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wdata6(.PAD(mem_wdata[6]), .A(mem_wdata_w[6]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wdata7(.PAD(mem_wdata[7]), .A(mem_wdata_w[7]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wdata8(.PAD(mem_wdata[8]), .A(mem_wdata_w[8]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wdata9(.PAD(mem_wdata[9]), .A(mem_wdata_w[9]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wdata10(.PAD(mem_wdata[10]), .A(mem_wdata_w[10]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wdata11(.PAD(mem_wdata[11]), .A(mem_wdata_w[11]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wdata12(.PAD(mem_wdata[12]), .A(mem_wdata_w[12]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wdata13(.PAD(mem_wdata[13]), .A(mem_wdata_w[13]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wdata14(.PAD(mem_wdata[14]), .A(mem_wdata_w[14]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wdata15(.PAD(mem_wdata[15]), .A(mem_wdata_w[15]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wdata16(.PAD(mem_wdata[16]), .A(mem_wdata_w[16]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wdata17(.PAD(mem_wdata[17]), .A(mem_wdata_w[17]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wdata18(.PAD(mem_wdata[18]), .A(mem_wdata_w[18]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wdata19(.PAD(mem_wdata[19]), .A(mem_wdata_w[19]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wdata20(.PAD(mem_wdata[20]), .A(mem_wdata_w[20]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wdata21(.PAD(mem_wdata[21]), .A(mem_wdata_w[21]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wdata22(.PAD(mem_wdata[22]), .A(mem_wdata_w[22]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wdata23(.PAD(mem_wdata[23]), .A(mem_wdata_w[23]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wdata24(.PAD(mem_wdata[24]), .A(mem_wdata_w[24]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wdata25(.PAD(mem_wdata[25]), .A(mem_wdata_w[25]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wdata26(.PAD(mem_wdata[26]), .A(mem_wdata_w[26]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wdata27(.PAD(mem_wdata[27]), .A(mem_wdata_w[27]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wdata28(.PAD(mem_wdata[28]), .A(mem_wdata_w[28]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wdata29(.PAD(mem_wdata[29]), .A(mem_wdata_w[29]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wdata30(.PAD(mem_wdata[30]), .A(mem_wdata_w[30]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wdata31(.PAD(mem_wdata[31]), .A(mem_wdata_w[31]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_addr0(.PAD(mem_la_addr[0]), .A(mem_la_addr_w[0]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_addr1(.PAD(mem_la_addr[1]), .A(mem_la_addr_w[1]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_addr2(.PAD(mem_la_addr[2]), .A(mem_la_addr_w[2]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_addr3(.PAD(mem_la_addr[3]), .A(mem_la_addr_w[3]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_addr4(.PAD(mem_la_addr[4]), .A(mem_la_addr_w[4]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_addr5(.PAD(mem_la_addr[5]), .A(mem_la_addr_w[5]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_addr6(.PAD(mem_la_addr[6]), .A(mem_la_addr_w[6]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_addr7(.PAD(mem_la_addr[7]), .A(mem_la_addr_w[7]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_addr8(.PAD(mem_la_addr[8]), .A(mem_la_addr_w[8]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_addr9(.PAD(mem_la_addr[9]), .A(mem_la_addr_w[9]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_addr10(.PAD(mem_la_addr[10]), .A(mem_la_addr_w[10]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_addr11(.PAD(mem_la_addr[11]), .A(mem_la_addr_w[11]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_addr12(.PAD(mem_la_addr[12]), .A(mem_la_addr_w[12]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_addr13(.PAD(mem_la_addr[13]), .A(mem_la_addr_w[13]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_addr14(.PAD(mem_la_addr[14]), .A(mem_la_addr_w[14]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_addr15(.PAD(mem_la_addr[15]), .A(mem_la_addr_w[15]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_addr16(.PAD(mem_la_addr[16]), .A(mem_la_addr_w[16]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_addr17(.PAD(mem_la_addr[17]), .A(mem_la_addr_w[17]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_addr18(.PAD(mem_la_addr[18]), .A(mem_la_addr_w[18]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_addr19(.PAD(mem_la_addr[19]), .A(mem_la_addr_w[19]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_addr20(.PAD(mem_la_addr[20]), .A(mem_la_addr_w[20]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_addr21(.PAD(mem_la_addr[21]), .A(mem_la_addr_w[21]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_addr22(.PAD(mem_la_addr[22]), .A(mem_la_addr_w[22]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_addr23(.PAD(mem_la_addr[23]), .A(mem_la_addr_w[23]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_addr24(.PAD(mem_la_addr[24]), .A(mem_la_addr_w[24]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_addr25(.PAD(mem_la_addr[25]), .A(mem_la_addr_w[25]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_addr26(.PAD(mem_la_addr[26]), .A(mem_la_addr_w[26]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_addr27(.PAD(mem_la_addr[27]), .A(mem_la_addr_w[27]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_addr28(.PAD(mem_la_addr[28]), .A(mem_la_addr_w[28]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_addr29(.PAD(mem_la_addr[29]), .A(mem_la_addr_w[29]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_addr30(.PAD(mem_la_addr[30]), .A(mem_la_addr_w[30]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_addr31(.PAD(mem_la_addr[31]), .A(mem_la_addr_w[31]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wdata0(.PAD(mem_la_wdata[0]), .A(mem_la_wdata_w[0]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wdata1(.PAD(mem_la_wdata[1]), .A(mem_la_wdata_w[1]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wdata2(.PAD(mem_la_wdata[2]), .A(mem_la_wdata_w[2]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wdata3(.PAD(mem_la_wdata[3]), .A(mem_la_wdata_w[3]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wdata4(.PAD(mem_la_wdata[4]), .A(mem_la_wdata_w[4]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wdata5(.PAD(mem_la_wdata[5]), .A(mem_la_wdata_w[5]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wdata6(.PAD(mem_la_wdata[6]), .A(mem_la_wdata_w[6]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wdata7(.PAD(mem_la_wdata[7]), .A(mem_la_wdata_w[7]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wdata8(.PAD(mem_la_wdata[8]), .A(mem_la_wdata_w[8]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wdata9(.PAD(mem_la_wdata[9]), .A(mem_la_wdata_w[9]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wdata10(.PAD(mem_la_wdata[10]), .A(mem_la_wdata_w[10]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wdata11(.PAD(mem_la_wdata[11]), .A(mem_la_wdata_w[11]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wdata12(.PAD(mem_la_wdata[12]), .A(mem_la_wdata_w[12]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wdata13(.PAD(mem_la_wdata[13]), .A(mem_la_wdata_w[13]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wdata14(.PAD(mem_la_wdata[14]), .A(mem_la_wdata_w[14]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wdata15(.PAD(mem_la_wdata[15]), .A(mem_la_wdata_w[15]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wdata16(.PAD(mem_la_wdata[16]), .A(mem_la_wdata_w[16]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wdata17(.PAD(mem_la_wdata[17]), .A(mem_la_wdata_w[17]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wdata18(.PAD(mem_la_wdata[18]), .A(mem_la_wdata_w[18]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wdata19(.PAD(mem_la_wdata[19]), .A(mem_la_wdata_w[19]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wdata20(.PAD(mem_la_wdata[20]), .A(mem_la_wdata_w[20]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wdata21(.PAD(mem_la_wdata[21]), .A(mem_la_wdata_w[21]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wdata22(.PAD(mem_la_wdata[22]), .A(mem_la_wdata_w[22]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wdata23(.PAD(mem_la_wdata[23]), .A(mem_la_wdata_w[23]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wdata24(.PAD(mem_la_wdata[24]), .A(mem_la_wdata_w[24]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wdata25(.PAD(mem_la_wdata[25]), .A(mem_la_wdata_w[25]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wdata26(.PAD(mem_la_wdata[26]), .A(mem_la_wdata_w[26]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wdata27(.PAD(mem_la_wdata[27]), .A(mem_la_wdata_w[27]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wdata28(.PAD(mem_la_wdata[28]), .A(mem_la_wdata_w[28]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wdata29(.PAD(mem_la_wdata[29]), .A(mem_la_wdata_w[29]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wdata30(.PAD(mem_la_wdata[30]), .A(mem_la_wdata_w[30]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wdata31(.PAD(mem_la_wdata[31]), .A(mem_la_wdata_w[31]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_insn0(.PAD(pcpi_insn[0]), .A(pcpi_insn_w[0]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_insn1(.PAD(pcpi_insn[1]), .A(pcpi_insn_w[1]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_insn2(.PAD(pcpi_insn[2]), .A(pcpi_insn_w[2]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_insn3(.PAD(pcpi_insn[3]), .A(pcpi_insn_w[3]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_insn4(.PAD(pcpi_insn[4]), .A(pcpi_insn_w[4]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_insn5(.PAD(pcpi_insn[5]), .A(pcpi_insn_w[5]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_insn6(.PAD(pcpi_insn[6]), .A(pcpi_insn_w[6]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_insn7(.PAD(pcpi_insn[7]), .A(pcpi_insn_w[7]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_insn8(.PAD(pcpi_insn[8]), .A(pcpi_insn_w[8]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_insn9(.PAD(pcpi_insn[9]), .A(pcpi_insn_w[9]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_insn10(.PAD(pcpi_insn[10]), .A(pcpi_insn_w[10]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_insn11(.PAD(pcpi_insn[11]), .A(pcpi_insn_w[11]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_insn12(.PAD(pcpi_insn[12]), .A(pcpi_insn_w[12]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_insn13(.PAD(pcpi_insn[13]), .A(pcpi_insn_w[13]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_insn14(.PAD(pcpi_insn[14]), .A(pcpi_insn_w[14]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_insn15(.PAD(pcpi_insn[15]), .A(pcpi_insn_w[15]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_insn16(.PAD(pcpi_insn[16]), .A(pcpi_insn_w[16]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_insn17(.PAD(pcpi_insn[17]), .A(pcpi_insn_w[17]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_insn18(.PAD(pcpi_insn[18]), .A(pcpi_insn_w[18]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_insn19(.PAD(pcpi_insn[19]), .A(pcpi_insn_w[19]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_insn20(.PAD(pcpi_insn[20]), .A(pcpi_insn_w[20]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_insn21(.PAD(pcpi_insn[21]), .A(pcpi_insn_w[21]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_insn22(.PAD(pcpi_insn[22]), .A(pcpi_insn_w[22]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_insn23(.PAD(pcpi_insn[23]), .A(pcpi_insn_w[23]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_insn24(.PAD(pcpi_insn[24]), .A(pcpi_insn_w[24]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_insn25(.PAD(pcpi_insn[25]), .A(pcpi_insn_w[25]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_insn26(.PAD(pcpi_insn[26]), .A(pcpi_insn_w[26]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_insn27(.PAD(pcpi_insn[27]), .A(pcpi_insn_w[27]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_insn28(.PAD(pcpi_insn[28]), .A(pcpi_insn_w[28]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_insn29(.PAD(pcpi_insn[29]), .A(pcpi_insn_w[29]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_insn30(.PAD(pcpi_insn[30]), .A(pcpi_insn_w[30]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_insn31(.PAD(pcpi_insn[31]), .A(pcpi_insn_w[31]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs10(.PAD(pcpi_rs1[0]), .A(pcpi_rs1_w[0]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs11(.PAD(pcpi_rs1[1]), .A(pcpi_rs1_w[1]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs12(.PAD(pcpi_rs1[2]), .A(pcpi_rs1_w[2]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs13(.PAD(pcpi_rs1[3]), .A(pcpi_rs1_w[3]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs14(.PAD(pcpi_rs1[4]), .A(pcpi_rs1_w[4]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs15(.PAD(pcpi_rs1[5]), .A(pcpi_rs1_w[5]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs16(.PAD(pcpi_rs1[6]), .A(pcpi_rs1_w[6]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs17(.PAD(pcpi_rs1[7]), .A(pcpi_rs1_w[7]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs18(.PAD(pcpi_rs1[8]), .A(pcpi_rs1_w[8]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs19(.PAD(pcpi_rs1[9]), .A(pcpi_rs1_w[9]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs110(.PAD(pcpi_rs1[10]), .A(pcpi_rs1_w[10]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs111(.PAD(pcpi_rs1[11]), .A(pcpi_rs1_w[11]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs112(.PAD(pcpi_rs1[12]), .A(pcpi_rs1_w[12]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs113(.PAD(pcpi_rs1[13]), .A(pcpi_rs1_w[13]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs114(.PAD(pcpi_rs1[14]), .A(pcpi_rs1_w[14]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs115(.PAD(pcpi_rs1[15]), .A(pcpi_rs1_w[15]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs116(.PAD(pcpi_rs1[16]), .A(pcpi_rs1_w[16]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs117(.PAD(pcpi_rs1[17]), .A(pcpi_rs1_w[17]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs118(.PAD(pcpi_rs1[18]), .A(pcpi_rs1_w[18]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs119(.PAD(pcpi_rs1[19]), .A(pcpi_rs1_w[19]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs120(.PAD(pcpi_rs1[20]), .A(pcpi_rs1_w[20]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs121(.PAD(pcpi_rs1[21]), .A(pcpi_rs1_w[21]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs122(.PAD(pcpi_rs1[22]), .A(pcpi_rs1_w[22]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs123(.PAD(pcpi_rs1[23]), .A(pcpi_rs1_w[23]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs124(.PAD(pcpi_rs1[24]), .A(pcpi_rs1_w[24]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs125(.PAD(pcpi_rs1[25]), .A(pcpi_rs1_w[25]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs126(.PAD(pcpi_rs1[26]), .A(pcpi_rs1_w[26]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs127(.PAD(pcpi_rs1[27]), .A(pcpi_rs1_w[27]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs128(.PAD(pcpi_rs1[28]), .A(pcpi_rs1_w[28]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs129(.PAD(pcpi_rs1[29]), .A(pcpi_rs1_w[29]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs130(.PAD(pcpi_rs1[30]), .A(pcpi_rs1_w[30]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs131(.PAD(pcpi_rs1[31]), .A(pcpi_rs1_w[31]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs20(.PAD(pcpi_rs2[0]), .A(pcpi_rs2_w[0]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs21(.PAD(pcpi_rs2[1]), .A(pcpi_rs2_w[1]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs22(.PAD(pcpi_rs2[2]), .A(pcpi_rs2_w[2]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs23(.PAD(pcpi_rs2[3]), .A(pcpi_rs2_w[3]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs24(.PAD(pcpi_rs2[4]), .A(pcpi_rs2_w[4]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs25(.PAD(pcpi_rs2[5]), .A(pcpi_rs2_w[5]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs26(.PAD(pcpi_rs2[6]), .A(pcpi_rs2_w[6]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs27(.PAD(pcpi_rs2[7]), .A(pcpi_rs2_w[7]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs28(.PAD(pcpi_rs2[8]), .A(pcpi_rs2_w[8]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs29(.PAD(pcpi_rs2[9]), .A(pcpi_rs2_w[9]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs210(.PAD(pcpi_rs2[10]), .A(pcpi_rs2_w[10]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs211(.PAD(pcpi_rs2[11]), .A(pcpi_rs2_w[11]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs212(.PAD(pcpi_rs2[12]), .A(pcpi_rs2_w[12]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs213(.PAD(pcpi_rs2[13]), .A(pcpi_rs2_w[13]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs214(.PAD(pcpi_rs2[14]), .A(pcpi_rs2_w[14]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs215(.PAD(pcpi_rs2[15]), .A(pcpi_rs2_w[15]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs216(.PAD(pcpi_rs2[16]), .A(pcpi_rs2_w[16]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs217(.PAD(pcpi_rs2[17]), .A(pcpi_rs2_w[17]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs218(.PAD(pcpi_rs2[18]), .A(pcpi_rs2_w[18]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs219(.PAD(pcpi_rs2[19]), .A(pcpi_rs2_w[19]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs220(.PAD(pcpi_rs2[20]), .A(pcpi_rs2_w[20]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs221(.PAD(pcpi_rs2[21]), .A(pcpi_rs2_w[21]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs222(.PAD(pcpi_rs2[22]), .A(pcpi_rs2_w[22]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs223(.PAD(pcpi_rs2[23]), .A(pcpi_rs2_w[23]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs224(.PAD(pcpi_rs2[24]), .A(pcpi_rs2_w[24]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs225(.PAD(pcpi_rs2[25]), .A(pcpi_rs2_w[25]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs226(.PAD(pcpi_rs2[26]), .A(pcpi_rs2_w[26]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs227(.PAD(pcpi_rs2[27]), .A(pcpi_rs2_w[27]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs228(.PAD(pcpi_rs2[28]), .A(pcpi_rs2_w[28]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs229(.PAD(pcpi_rs2[29]), .A(pcpi_rs2_w[29]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs230(.PAD(pcpi_rs2[30]), .A(pcpi_rs2_w[30]), .VDD(VDD), .VSS(VSS));
PADDO pad_pcpi_rs231(.PAD(pcpi_rs2[31]), .A(pcpi_rs2_w[31]), .VDD(VDD), .VSS(VSS));
PADDO pad_eoi0(.PAD(eoi[0]), .A(eoi_w[0]), .VDD(VDD), .VSS(VSS));
PADDO pad_eoi1(.PAD(eoi[1]), .A(eoi_w[1]), .VDD(VDD), .VSS(VSS));
PADDO pad_eoi2(.PAD(eoi[2]), .A(eoi_w[2]), .VDD(VDD), .VSS(VSS));
PADDO pad_eoi3(.PAD(eoi[3]), .A(eoi_w[3]), .VDD(VDD), .VSS(VSS));
PADDO pad_eoi4(.PAD(eoi[4]), .A(eoi_w[4]), .VDD(VDD), .VSS(VSS));
PADDO pad_eoi5(.PAD(eoi[5]), .A(eoi_w[5]), .VDD(VDD), .VSS(VSS));
PADDO pad_eoi6(.PAD(eoi[6]), .A(eoi_w[6]), .VDD(VDD), .VSS(VSS));
PADDO pad_eoi7(.PAD(eoi[7]), .A(eoi_w[7]), .VDD(VDD), .VSS(VSS));
PADDO pad_eoi8(.PAD(eoi[8]), .A(eoi_w[8]), .VDD(VDD), .VSS(VSS));
PADDO pad_eoi9(.PAD(eoi[9]), .A(eoi_w[9]), .VDD(VDD), .VSS(VSS));
PADDO pad_eoi10(.PAD(eoi[10]), .A(eoi_w[10]), .VDD(VDD), .VSS(VSS));
PADDO pad_eoi11(.PAD(eoi[11]), .A(eoi_w[11]), .VDD(VDD), .VSS(VSS));
PADDO pad_eoi12(.PAD(eoi[12]), .A(eoi_w[12]), .VDD(VDD), .VSS(VSS));
PADDO pad_eoi13(.PAD(eoi[13]), .A(eoi_w[13]), .VDD(VDD), .VSS(VSS));
PADDO pad_eoi14(.PAD(eoi[14]), .A(eoi_w[14]), .VDD(VDD), .VSS(VSS));
PADDO pad_eoi15(.PAD(eoi[15]), .A(eoi_w[15]), .VDD(VDD), .VSS(VSS));
PADDO pad_eoi16(.PAD(eoi[16]), .A(eoi_w[16]), .VDD(VDD), .VSS(VSS));
PADDO pad_eoi17(.PAD(eoi[17]), .A(eoi_w[17]), .VDD(VDD), .VSS(VSS));
PADDO pad_eoi18(.PAD(eoi[18]), .A(eoi_w[18]), .VDD(VDD), .VSS(VSS));
PADDO pad_eoi19(.PAD(eoi[19]), .A(eoi_w[19]), .VDD(VDD), .VSS(VSS));
PADDO pad_eoi20(.PAD(eoi[20]), .A(eoi_w[20]), .VDD(VDD), .VSS(VSS));
PADDO pad_eoi21(.PAD(eoi[21]), .A(eoi_w[21]), .VDD(VDD), .VSS(VSS));
PADDO pad_eoi22(.PAD(eoi[22]), .A(eoi_w[22]), .VDD(VDD), .VSS(VSS));
PADDO pad_eoi23(.PAD(eoi[23]), .A(eoi_w[23]), .VDD(VDD), .VSS(VSS));
PADDO pad_eoi24(.PAD(eoi[24]), .A(eoi_w[24]), .VDD(VDD), .VSS(VSS));
PADDO pad_eoi25(.PAD(eoi[25]), .A(eoi_w[25]), .VDD(VDD), .VSS(VSS));
PADDO pad_eoi26(.PAD(eoi[26]), .A(eoi_w[26]), .VDD(VDD), .VSS(VSS));
PADDO pad_eoi27(.PAD(eoi[27]), .A(eoi_w[27]), .VDD(VDD), .VSS(VSS));
PADDO pad_eoi28(.PAD(eoi[28]), .A(eoi_w[28]), .VDD(VDD), .VSS(VSS));
PADDO pad_eoi29(.PAD(eoi[29]), .A(eoi_w[29]), .VDD(VDD), .VSS(VSS));
PADDO pad_eoi30(.PAD(eoi[30]), .A(eoi_w[30]), .VDD(VDD), .VSS(VSS));
PADDO pad_eoi31(.PAD(eoi[31]), .A(eoi_w[31]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wstrb0(.PAD(mem_wstrb[0]), .A(mem_wstrb_w[0]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wstrb1(.PAD(mem_wstrb[1]), .A(mem_wstrb_w[1]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wstrb2(.PAD(mem_wstrb[2]), .A(mem_wstrb_w[2]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_wstrb3(.PAD(mem_wstrb[3]), .A(mem_wstrb_w[3]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wstrb0(.PAD(mem_la_wstrb[0]), .A(mem_la_wstrb_w[0]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wstrb1(.PAD(mem_la_wstrb[1]), .A(mem_la_wstrb_w[1]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wstrb2(.PAD(mem_la_wstrb[2]), .A(mem_la_wstrb_w[2]), .VDD(VDD), .VSS(VSS));
PADDO pad_mem_la_wstrb3(.PAD(mem_la_wstrb[3]), .A(mem_la_wstrb_w[3]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data0(.PAD(trace_data[0]), .A(trace_data_w[0]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data1(.PAD(trace_data[1]), .A(trace_data_w[1]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data2(.PAD(trace_data[2]), .A(trace_data_w[2]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data3(.PAD(trace_data[3]), .A(trace_data_w[3]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data4(.PAD(trace_data[4]), .A(trace_data_w[4]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data5(.PAD(trace_data[5]), .A(trace_data_w[5]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data6(.PAD(trace_data[6]), .A(trace_data_w[6]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data7(.PAD(trace_data[7]), .A(trace_data_w[7]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data8(.PAD(trace_data[8]), .A(trace_data_w[8]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data9(.PAD(trace_data[9]), .A(trace_data_w[9]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data10(.PAD(trace_data[10]), .A(trace_data_w[10]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data11(.PAD(trace_data[11]), .A(trace_data_w[11]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data12(.PAD(trace_data[12]), .A(trace_data_w[12]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data13(.PAD(trace_data[13]), .A(trace_data_w[13]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data14(.PAD(trace_data[14]), .A(trace_data_w[14]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data15(.PAD(trace_data[15]), .A(trace_data_w[15]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data16(.PAD(trace_data[16]), .A(trace_data_w[16]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data17(.PAD(trace_data[17]), .A(trace_data_w[17]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data18(.PAD(trace_data[18]), .A(trace_data_w[18]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data19(.PAD(trace_data[19]), .A(trace_data_w[19]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data20(.PAD(trace_data[20]), .A(trace_data_w[20]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data21(.PAD(trace_data[21]), .A(trace_data_w[21]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data22(.PAD(trace_data[22]), .A(trace_data_w[22]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data23(.PAD(trace_data[23]), .A(trace_data_w[23]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data24(.PAD(trace_data[24]), .A(trace_data_w[24]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data25(.PAD(trace_data[25]), .A(trace_data_w[25]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data26(.PAD(trace_data[26]), .A(trace_data_w[26]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data27(.PAD(trace_data[27]), .A(trace_data_w[27]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data28(.PAD(trace_data[28]), .A(trace_data_w[28]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data29(.PAD(trace_data[29]), .A(trace_data_w[29]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data30(.PAD(trace_data[30]), .A(trace_data_w[30]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data31(.PAD(trace_data[31]), .A(trace_data_w[31]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data32(.PAD(trace_data[32]), .A(trace_data_w[32]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data33(.PAD(trace_data[33]), .A(trace_data_w[33]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data34(.PAD(trace_data[34]), .A(trace_data_w[34]), .VDD(VDD), .VSS(VSS));
PADDO pad_trace_data35(.PAD(trace_data[35]), .A(trace_data_w[35]), .VDD(VDD), .VSS(VSS));

//Insert Corners
  padIORINGCORNER pad_corner0();
  padIORINGCORNER pad_corner1();
  padIORINGCORNER pad_corner2();
  padIORINGCORNER pad_corner3();

endmodule


module picorv32(clk, resetn, trap, mem_valid, mem_instr, mem_ready,
     mem_addr, mem_wdata, mem_wstrb, mem_rdata, mem_la_read,
     mem_la_write, mem_la_addr, mem_la_wdata, mem_la_wstrb, pcpi_valid,
     pcpi_insn, pcpi_rs1, pcpi_rs2, pcpi_wr, pcpi_rd, pcpi_wait,
     pcpi_ready, irq, eoi, trace_valid, trace_data);
  input clk, resetn, mem_ready, pcpi_wr, pcpi_wait, pcpi_ready;
  input [31:0] mem_rdata, pcpi_rd, irq;
  output trap, mem_valid, mem_instr, mem_la_read, mem_la_write,
       pcpi_valid, trace_valid;
  output [31:0] mem_addr, mem_wdata, mem_la_addr, mem_la_wdata,
       pcpi_insn, pcpi_rs1, pcpi_rs2, eoi;
  output [3:0] mem_wstrb, mem_la_wstrb;
  output [35:0] trace_data;
  wire clk, resetn, mem_ready, pcpi_wr, pcpi_wait, pcpi_ready;
  wire [31:0] mem_rdata, pcpi_rd, irq;
  wire trap, mem_valid, mem_instr, mem_la_read, mem_la_write,
       pcpi_valid, trace_valid;
  wire [31:0] mem_addr, mem_wdata, mem_la_addr, mem_la_wdata,
       pcpi_insn, pcpi_rs1, pcpi_rs2, eoi;
  wire [3:0] mem_wstrb, mem_la_wstrb;
  wire [35:0] trace_data;
  wire [31:0] \genblk2.pcpi_div_dividend ;
  wire [31:0] \genblk2.pcpi_div_quotient ;
  wire [31:0] alu_out_q;
  wire [63:0] \genblk1.pcpi_mul_rd ;
  wire [31:0] pcpi_div_rd;
  wire [31:0] reg_out;
  wire [31:0] current_pc;
  wire [7:0] cpu_state;
  wire [31:0] decoded_imm;
  wire [31:0] reg_op1;
  wire [62:0] \genblk2.pcpi_div_divisor ;
  wire [31:0] mem_rdata_latched;
  wire [15:0] mem_16bit_buffer;
  wire [31:0] mem_rdata_q;
  wire [31:0] reg_next_pc;
  wire [3:0] pcpi_timeout_counter;
  wire [63:0] count_instr;
  wire [63:0] count_cycle;
  wire [31:0] decoded_imm_j;
  wire [1:0] mem_state;
  wire [1:0] mem_wordsize;
  wire [31:0] \cpuregs[1] ;
  wire [31:0] \cpuregs[2] ;
  wire [31:0] \cpuregs[3] ;
  wire [31:0] \cpuregs[4] ;
  wire [31:0] \cpuregs[5] ;
  wire [31:0] \cpuregs[6] ;
  wire [31:0] \cpuregs[7] ;
  wire [31:0] \cpuregs[8] ;
  wire [31:0] \cpuregs[9] ;
  wire [31:0] \cpuregs[10] ;
  wire [31:0] \cpuregs[11] ;
  wire [31:0] \cpuregs[12] ;
  wire [31:0] \cpuregs[13] ;
  wire [31:0] \cpuregs[14] ;
  wire [31:0] \cpuregs[15] ;
  wire [31:0] \cpuregs[16] ;
  wire [31:0] \cpuregs[17] ;
  wire [31:0] \cpuregs[18] ;
  wire [31:0] \cpuregs[19] ;
  wire [31:0] \cpuregs[20] ;
  wire [31:0] \cpuregs[21] ;
  wire [31:0] \cpuregs[22] ;
  wire [31:0] \cpuregs[23] ;
  wire [31:0] \cpuregs[24] ;
  wire [31:0] \cpuregs[25] ;
  wire [31:0] \cpuregs[26] ;
  wire [31:0] \cpuregs[27] ;
  wire [31:0] \cpuregs[28] ;
  wire [31:0] \cpuregs[29] ;
  wire [31:0] \cpuregs[30] ;
  wire [31:0] \cpuregs[31] ;
  wire [4:0] decoded_rd;
  wire [4:0] decoded_rs1;
  wire [4:0] decoded_rs2;
  wire [3:0] \genblk1.pcpi_mul_active ;
  wire [32:0] \genblk1.pcpi_mul_rs1 ;
  wire [32:0] \genblk1.pcpi_mul_rs2 ;
  wire [31:0] \genblk2.pcpi_div_quotient_msk ;
  wire [4:0] latched_rd;
  wire [31:0] reg_pc;
  wire [4:0] reg_sh;
  wire UNCONNECTED, add_1312_30_n_102, add_1312_30_n_851,
       add_1312_30_n_856, add_1312_30_n_861, add_1312_30_n_866,
       add_1312_30_n_871, add_1312_30_n_876;
  wire add_1312_30_n_881, add_1312_30_n_886, add_1312_30_n_891,
       add_1312_30_n_896, add_1312_30_n_901, add_1312_30_n_906,
       add_1312_30_n_911, add_1312_30_n_916;
  wire add_1312_30_n_921, add_1312_30_n_926, add_1312_30_n_931,
       add_1312_30_n_936, add_1312_30_n_941, add_1312_30_n_946,
       add_1312_30_n_951, add_1312_30_n_956;
  wire add_1312_30_n_961, add_1312_30_n_966, add_1312_30_n_971,
       add_1312_30_n_976, add_1312_30_n_981, add_1312_30_n_986,
       add_1312_30_n_991, add_1312_30_n_1020;
  wire add_1564_33_Y_add_1555_32_n_585,
       add_1564_33_Y_add_1555_32_n_587,
       add_1564_33_Y_add_1555_32_n_590,
       add_1564_33_Y_add_1555_32_n_592,
       add_1564_33_Y_add_1555_32_n_594,
       add_1564_33_Y_add_1555_32_n_596,
       add_1564_33_Y_add_1555_32_n_598, add_1564_33_Y_add_1555_32_n_600;
  wire add_1564_33_Y_add_1555_32_n_602,
       add_1564_33_Y_add_1555_32_n_604,
       add_1564_33_Y_add_1555_32_n_606,
       add_1564_33_Y_add_1555_32_n_608,
       add_1564_33_Y_add_1555_32_n_610,
       add_1564_33_Y_add_1555_32_n_612,
       add_1564_33_Y_add_1555_32_n_614, add_1564_33_Y_add_1555_32_n_616;
  wire add_1564_33_Y_add_1555_32_n_618,
       add_1564_33_Y_add_1555_32_n_620,
       add_1564_33_Y_add_1555_32_n_622,
       add_1564_33_Y_add_1555_32_n_624,
       add_1564_33_Y_add_1555_32_n_626,
       add_1564_33_Y_add_1555_32_n_628,
       add_1564_33_Y_add_1555_32_n_630, add_1564_33_Y_add_1555_32_n_632;
  wire add_1564_33_Y_add_1555_32_n_634,
       add_1564_33_Y_add_1555_32_n_636,
       add_1564_33_Y_add_1555_32_n_638,
       add_1564_33_Y_add_1555_32_n_640,
       add_1564_33_Y_add_1555_32_n_642,
       add_1564_33_Y_add_1555_32_n_645,
       add_1564_33_Y_add_1555_32_n_646, add_1801_23_n_1105;
  wire add_1801_23_n_1107, add_1801_23_n_1109, add_1801_23_n_1111,
       add_1801_23_n_1113, add_1801_23_n_1115, add_1801_23_n_1117,
       add_1801_23_n_1119, add_1801_23_n_1121;
  wire add_1801_23_n_1123, add_1801_23_n_1125, add_1801_23_n_1127,
       add_1801_23_n_1129, add_1801_23_n_1131, add_1801_23_n_1133,
       add_1801_23_n_1135, add_1801_23_n_1137;
  wire add_1801_23_n_1139, add_1801_23_n_1141, add_1801_23_n_1143,
       add_1801_23_n_1145, add_1801_23_n_1147, add_1801_23_n_1149,
       add_1801_23_n_1151, add_1801_23_n_1153;
  wire add_1801_23_n_1155, add_1801_23_n_1157, add_1801_23_n_1159,
       add_1801_23_n_1161, add_1801_23_n_1164, add_1801_23_n_1165,
       add_1864_26_n_596, add_1864_26_n_598;
  wire add_1864_26_n_600, add_1864_26_n_602, add_1864_26_n_604,
       add_1864_26_n_606, add_1864_26_n_608, add_1864_26_n_610,
       add_1864_26_n_612, add_1864_26_n_614;
  wire add_1864_26_n_616, add_1864_26_n_618, add_1864_26_n_620,
       add_1864_26_n_622, add_1864_26_n_624, add_1864_26_n_626,
       add_1864_26_n_628, add_1864_26_n_630;
  wire add_1864_26_n_632, add_1864_26_n_634, add_1864_26_n_636,
       add_1864_26_n_638, add_1864_26_n_640, add_1864_26_n_642,
       add_1864_26_n_644, add_1864_26_n_646;
  wire add_1864_26_n_648, add_1864_26_n_650, add_1864_26_n_652,
       add_1864_26_n_654, add_1864_26_n_657, add_1864_26_n_658,
       clear_prefetched_high_word_q, compressed_instr;
  wire decoder_pseudo_trigger, decoder_trigger,
       \genblk1.pcpi_mul_mul_2366_47_n_0 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2 ,
       \genblk1.pcpi_mul_mul_2366_47_n_3 ,
       \genblk1.pcpi_mul_mul_2366_47_n_4 ,
       \genblk1.pcpi_mul_mul_2366_47_n_5 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_6 ,
       \genblk1.pcpi_mul_mul_2366_47_n_7 ,
       \genblk1.pcpi_mul_mul_2366_47_n_8 ,
       \genblk1.pcpi_mul_mul_2366_47_n_9 ,
       \genblk1.pcpi_mul_mul_2366_47_n_10 ,
       \genblk1.pcpi_mul_mul_2366_47_n_11 ,
       \genblk1.pcpi_mul_mul_2366_47_n_12 ,
       \genblk1.pcpi_mul_mul_2366_47_n_13 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_14 ,
       \genblk1.pcpi_mul_mul_2366_47_n_16 ,
       \genblk1.pcpi_mul_mul_2366_47_n_18 ,
       \genblk1.pcpi_mul_mul_2366_47_n_20 ,
       \genblk1.pcpi_mul_mul_2366_47_n_22 ,
       \genblk1.pcpi_mul_mul_2366_47_n_24 ,
       \genblk1.pcpi_mul_mul_2366_47_n_35 ,
       \genblk1.pcpi_mul_mul_2366_47_n_37 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_39 ,
       \genblk1.pcpi_mul_mul_2366_47_n_41 ,
       \genblk1.pcpi_mul_mul_2366_47_n_43 ,
       \genblk1.pcpi_mul_mul_2366_47_n_45 ,
       \genblk1.pcpi_mul_mul_2366_47_n_47 ,
       \genblk1.pcpi_mul_mul_2366_47_n_49 ,
       \genblk1.pcpi_mul_mul_2366_47_n_51 ,
       \genblk1.pcpi_mul_mul_2366_47_n_53 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_55 ,
       \genblk1.pcpi_mul_mul_2366_47_n_57 ,
       \genblk1.pcpi_mul_mul_2366_47_n_59 ,
       \genblk1.pcpi_mul_mul_2366_47_n_61 ,
       \genblk1.pcpi_mul_mul_2366_47_n_63 ,
       \genblk1.pcpi_mul_mul_2366_47_n_65 ,
       \genblk1.pcpi_mul_mul_2366_47_n_67 ,
       \genblk1.pcpi_mul_mul_2366_47_n_69 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_71 ,
       \genblk1.pcpi_mul_mul_2366_47_n_73 ,
       \genblk1.pcpi_mul_mul_2366_47_n_75 ,
       \genblk1.pcpi_mul_mul_2366_47_n_77 ,
       \genblk1.pcpi_mul_mul_2366_47_n_79 ,
       \genblk1.pcpi_mul_mul_2366_47_n_81 ,
       \genblk1.pcpi_mul_mul_2366_47_n_83 ,
       \genblk1.pcpi_mul_mul_2366_47_n_85 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_87 ,
       \genblk1.pcpi_mul_mul_2366_47_n_89 ,
       \genblk1.pcpi_mul_mul_2366_47_n_91 ,
       \genblk1.pcpi_mul_mul_2366_47_n_93 ,
       \genblk1.pcpi_mul_mul_2366_47_n_95 ,
       \genblk1.pcpi_mul_mul_2366_47_n_97 ,
       \genblk1.pcpi_mul_mul_2366_47_n_99 ,
       \genblk1.pcpi_mul_mul_2366_47_n_101 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_137 ,
       \genblk1.pcpi_mul_mul_2366_47_n_147 ,
       \genblk1.pcpi_mul_mul_2366_47_n_148 ,
       \genblk1.pcpi_mul_mul_2366_47_n_149 ,
       \genblk1.pcpi_mul_mul_2366_47_n_150 ,
       \genblk1.pcpi_mul_mul_2366_47_n_151 ,
       \genblk1.pcpi_mul_mul_2366_47_n_152 ,
       \genblk1.pcpi_mul_mul_2366_47_n_153 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_154 ,
       \genblk1.pcpi_mul_mul_2366_47_n_155 ,
       \genblk1.pcpi_mul_mul_2366_47_n_156 ,
       \genblk1.pcpi_mul_mul_2366_47_n_157 ,
       \genblk1.pcpi_mul_mul_2366_47_n_158 ,
       \genblk1.pcpi_mul_mul_2366_47_n_159 ,
       \genblk1.pcpi_mul_mul_2366_47_n_160 ,
       \genblk1.pcpi_mul_mul_2366_47_n_161 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_162 ,
       \genblk1.pcpi_mul_mul_2366_47_n_163 ,
       \genblk1.pcpi_mul_mul_2366_47_n_164 ,
       \genblk1.pcpi_mul_mul_2366_47_n_165 ,
       \genblk1.pcpi_mul_mul_2366_47_n_166 ,
       \genblk1.pcpi_mul_mul_2366_47_n_167 ,
       \genblk1.pcpi_mul_mul_2366_47_n_168 ,
       \genblk1.pcpi_mul_mul_2366_47_n_169 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_170 ,
       \genblk1.pcpi_mul_mul_2366_47_n_171 ,
       \genblk1.pcpi_mul_mul_2366_47_n_172 ,
       \genblk1.pcpi_mul_mul_2366_47_n_193 ,
       \genblk1.pcpi_mul_mul_2366_47_n_194 ,
       \genblk1.pcpi_mul_mul_2366_47_n_195 ,
       \genblk1.pcpi_mul_mul_2366_47_n_196 ,
       \genblk1.pcpi_mul_mul_2366_47_n_197 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_198 ,
       \genblk1.pcpi_mul_mul_2366_47_n_199 ,
       \genblk1.pcpi_mul_mul_2366_47_n_221 ,
       \genblk1.pcpi_mul_mul_2366_47_n_223 ,
       \genblk1.pcpi_mul_mul_2366_47_n_224 ,
       \genblk1.pcpi_mul_mul_2366_47_n_226 ,
       \genblk1.pcpi_mul_mul_2366_47_n_227 ,
       \genblk1.pcpi_mul_mul_2366_47_n_228 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_236 ,
       \genblk1.pcpi_mul_mul_2366_47_n_237 ,
       \genblk1.pcpi_mul_mul_2366_47_n_238 ,
       \genblk1.pcpi_mul_mul_2366_47_n_239 ,
       \genblk1.pcpi_mul_mul_2366_47_n_240 ,
       \genblk1.pcpi_mul_mul_2366_47_n_241 ,
       \genblk1.pcpi_mul_mul_2366_47_n_242 ,
       \genblk1.pcpi_mul_mul_2366_47_n_243 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_244 ,
       \genblk1.pcpi_mul_mul_2366_47_n_245 ,
       \genblk1.pcpi_mul_mul_2366_47_n_246 ,
       \genblk1.pcpi_mul_mul_2366_47_n_247 ,
       \genblk1.pcpi_mul_mul_2366_47_n_248 ,
       \genblk1.pcpi_mul_mul_2366_47_n_249 ,
       \genblk1.pcpi_mul_mul_2366_47_n_250 ,
       \genblk1.pcpi_mul_mul_2366_47_n_251 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_252 ,
       \genblk1.pcpi_mul_mul_2366_47_n_253 ,
       \genblk1.pcpi_mul_mul_2366_47_n_254 ,
       \genblk1.pcpi_mul_mul_2366_47_n_255 ,
       \genblk1.pcpi_mul_mul_2366_47_n_256 ,
       \genblk1.pcpi_mul_mul_2366_47_n_257 ,
       \genblk1.pcpi_mul_mul_2366_47_n_258 ,
       \genblk1.pcpi_mul_mul_2366_47_n_259 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_260 ,
       \genblk1.pcpi_mul_mul_2366_47_n_261 ,
       \genblk1.pcpi_mul_mul_2366_47_n_262 ,
       \genblk1.pcpi_mul_mul_2366_47_n_263 ,
       \genblk1.pcpi_mul_mul_2366_47_n_264 ,
       \genblk1.pcpi_mul_mul_2366_47_n_265 ,
       \genblk1.pcpi_mul_mul_2366_47_n_266 ,
       \genblk1.pcpi_mul_mul_2366_47_n_267 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_268 ,
       \genblk1.pcpi_mul_mul_2366_47_n_269 ,
       \genblk1.pcpi_mul_mul_2366_47_n_270 ,
       \genblk1.pcpi_mul_mul_2366_47_n_271 ,
       \genblk1.pcpi_mul_mul_2366_47_n_272 ,
       \genblk1.pcpi_mul_mul_2366_47_n_273 ,
       \genblk1.pcpi_mul_mul_2366_47_n_274 ,
       \genblk1.pcpi_mul_mul_2366_47_n_275 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_276 ,
       \genblk1.pcpi_mul_mul_2366_47_n_277 ,
       \genblk1.pcpi_mul_mul_2366_47_n_278 ,
       \genblk1.pcpi_mul_mul_2366_47_n_279 ,
       \genblk1.pcpi_mul_mul_2366_47_n_280 ,
       \genblk1.pcpi_mul_mul_2366_47_n_281 ,
       \genblk1.pcpi_mul_mul_2366_47_n_282 ,
       \genblk1.pcpi_mul_mul_2366_47_n_283 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_284 ,
       \genblk1.pcpi_mul_mul_2366_47_n_285 ,
       \genblk1.pcpi_mul_mul_2366_47_n_286 ,
       \genblk1.pcpi_mul_mul_2366_47_n_287 ,
       \genblk1.pcpi_mul_mul_2366_47_n_288 ,
       \genblk1.pcpi_mul_mul_2366_47_n_289 ,
       \genblk1.pcpi_mul_mul_2366_47_n_290 ,
       \genblk1.pcpi_mul_mul_2366_47_n_291 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_292 ,
       \genblk1.pcpi_mul_mul_2366_47_n_293 ,
       \genblk1.pcpi_mul_mul_2366_47_n_294 ,
       \genblk1.pcpi_mul_mul_2366_47_n_295 ,
       \genblk1.pcpi_mul_mul_2366_47_n_296 ,
       \genblk1.pcpi_mul_mul_2366_47_n_297 ,
       \genblk1.pcpi_mul_mul_2366_47_n_298 ,
       \genblk1.pcpi_mul_mul_2366_47_n_299 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_300 ,
       \genblk1.pcpi_mul_mul_2366_47_n_301 ,
       \genblk1.pcpi_mul_mul_2366_47_n_302 ,
       \genblk1.pcpi_mul_mul_2366_47_n_303 ,
       \genblk1.pcpi_mul_mul_2366_47_n_304 ,
       \genblk1.pcpi_mul_mul_2366_47_n_305 ,
       \genblk1.pcpi_mul_mul_2366_47_n_306 ,
       \genblk1.pcpi_mul_mul_2366_47_n_307 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_308 ,
       \genblk1.pcpi_mul_mul_2366_47_n_309 ,
       \genblk1.pcpi_mul_mul_2366_47_n_310 ,
       \genblk1.pcpi_mul_mul_2366_47_n_311 ,
       \genblk1.pcpi_mul_mul_2366_47_n_312 ,
       \genblk1.pcpi_mul_mul_2366_47_n_313 ,
       \genblk1.pcpi_mul_mul_2366_47_n_314 ,
       \genblk1.pcpi_mul_mul_2366_47_n_315 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_316 ,
       \genblk1.pcpi_mul_mul_2366_47_n_317 ,
       \genblk1.pcpi_mul_mul_2366_47_n_318 ,
       \genblk1.pcpi_mul_mul_2366_47_n_319 ,
       \genblk1.pcpi_mul_mul_2366_47_n_320 ,
       \genblk1.pcpi_mul_mul_2366_47_n_321 ,
       \genblk1.pcpi_mul_mul_2366_47_n_322 ,
       \genblk1.pcpi_mul_mul_2366_47_n_323 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_324 ,
       \genblk1.pcpi_mul_mul_2366_47_n_325 ,
       \genblk1.pcpi_mul_mul_2366_47_n_326 ,
       \genblk1.pcpi_mul_mul_2366_47_n_327 ,
       \genblk1.pcpi_mul_mul_2366_47_n_328 ,
       \genblk1.pcpi_mul_mul_2366_47_n_329 ,
       \genblk1.pcpi_mul_mul_2366_47_n_330 ,
       \genblk1.pcpi_mul_mul_2366_47_n_331 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_332 ,
       \genblk1.pcpi_mul_mul_2366_47_n_333 ,
       \genblk1.pcpi_mul_mul_2366_47_n_334 ,
       \genblk1.pcpi_mul_mul_2366_47_n_335 ,
       \genblk1.pcpi_mul_mul_2366_47_n_336 ,
       \genblk1.pcpi_mul_mul_2366_47_n_337 ,
       \genblk1.pcpi_mul_mul_2366_47_n_338 ,
       \genblk1.pcpi_mul_mul_2366_47_n_339 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_340 ,
       \genblk1.pcpi_mul_mul_2366_47_n_341 ,
       \genblk1.pcpi_mul_mul_2366_47_n_342 ,
       \genblk1.pcpi_mul_mul_2366_47_n_343 ,
       \genblk1.pcpi_mul_mul_2366_47_n_344 ,
       \genblk1.pcpi_mul_mul_2366_47_n_345 ,
       \genblk1.pcpi_mul_mul_2366_47_n_346 ,
       \genblk1.pcpi_mul_mul_2366_47_n_347 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_348 ,
       \genblk1.pcpi_mul_mul_2366_47_n_349 ,
       \genblk1.pcpi_mul_mul_2366_47_n_350 ,
       \genblk1.pcpi_mul_mul_2366_47_n_351 ,
       \genblk1.pcpi_mul_mul_2366_47_n_352 ,
       \genblk1.pcpi_mul_mul_2366_47_n_353 ,
       \genblk1.pcpi_mul_mul_2366_47_n_354 ,
       \genblk1.pcpi_mul_mul_2366_47_n_355 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_356 ,
       \genblk1.pcpi_mul_mul_2366_47_n_357 ,
       \genblk1.pcpi_mul_mul_2366_47_n_358 ,
       \genblk1.pcpi_mul_mul_2366_47_n_359 ,
       \genblk1.pcpi_mul_mul_2366_47_n_360 ,
       \genblk1.pcpi_mul_mul_2366_47_n_361 ,
       \genblk1.pcpi_mul_mul_2366_47_n_362 ,
       \genblk1.pcpi_mul_mul_2366_47_n_363 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_364 ,
       \genblk1.pcpi_mul_mul_2366_47_n_365 ,
       \genblk1.pcpi_mul_mul_2366_47_n_366 ,
       \genblk1.pcpi_mul_mul_2366_47_n_367 ,
       \genblk1.pcpi_mul_mul_2366_47_n_368 ,
       \genblk1.pcpi_mul_mul_2366_47_n_369 ,
       \genblk1.pcpi_mul_mul_2366_47_n_370 ,
       \genblk1.pcpi_mul_mul_2366_47_n_371 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_372 ,
       \genblk1.pcpi_mul_mul_2366_47_n_373 ,
       \genblk1.pcpi_mul_mul_2366_47_n_374 ,
       \genblk1.pcpi_mul_mul_2366_47_n_375 ,
       \genblk1.pcpi_mul_mul_2366_47_n_376 ,
       \genblk1.pcpi_mul_mul_2366_47_n_377 ,
       \genblk1.pcpi_mul_mul_2366_47_n_378 ,
       \genblk1.pcpi_mul_mul_2366_47_n_379 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_380 ,
       \genblk1.pcpi_mul_mul_2366_47_n_381 ,
       \genblk1.pcpi_mul_mul_2366_47_n_382 ,
       \genblk1.pcpi_mul_mul_2366_47_n_383 ,
       \genblk1.pcpi_mul_mul_2366_47_n_384 ,
       \genblk1.pcpi_mul_mul_2366_47_n_385 ,
       \genblk1.pcpi_mul_mul_2366_47_n_386 ,
       \genblk1.pcpi_mul_mul_2366_47_n_387 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_388 ,
       \genblk1.pcpi_mul_mul_2366_47_n_389 ,
       \genblk1.pcpi_mul_mul_2366_47_n_390 ,
       \genblk1.pcpi_mul_mul_2366_47_n_391 ,
       \genblk1.pcpi_mul_mul_2366_47_n_392 ,
       \genblk1.pcpi_mul_mul_2366_47_n_393 ,
       \genblk1.pcpi_mul_mul_2366_47_n_394 ,
       \genblk1.pcpi_mul_mul_2366_47_n_395 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_396 ,
       \genblk1.pcpi_mul_mul_2366_47_n_397 ,
       \genblk1.pcpi_mul_mul_2366_47_n_398 ,
       \genblk1.pcpi_mul_mul_2366_47_n_399 ,
       \genblk1.pcpi_mul_mul_2366_47_n_400 ,
       \genblk1.pcpi_mul_mul_2366_47_n_401 ,
       \genblk1.pcpi_mul_mul_2366_47_n_402 ,
       \genblk1.pcpi_mul_mul_2366_47_n_403 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_404 ,
       \genblk1.pcpi_mul_mul_2366_47_n_405 ,
       \genblk1.pcpi_mul_mul_2366_47_n_406 ,
       \genblk1.pcpi_mul_mul_2366_47_n_407 ,
       \genblk1.pcpi_mul_mul_2366_47_n_408 ,
       \genblk1.pcpi_mul_mul_2366_47_n_409 ,
       \genblk1.pcpi_mul_mul_2366_47_n_410 ,
       \genblk1.pcpi_mul_mul_2366_47_n_411 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_412 ,
       \genblk1.pcpi_mul_mul_2366_47_n_413 ,
       \genblk1.pcpi_mul_mul_2366_47_n_414 ,
       \genblk1.pcpi_mul_mul_2366_47_n_415 ,
       \genblk1.pcpi_mul_mul_2366_47_n_416 ,
       \genblk1.pcpi_mul_mul_2366_47_n_417 ,
       \genblk1.pcpi_mul_mul_2366_47_n_418 ,
       \genblk1.pcpi_mul_mul_2366_47_n_419 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_420 ,
       \genblk1.pcpi_mul_mul_2366_47_n_421 ,
       \genblk1.pcpi_mul_mul_2366_47_n_422 ,
       \genblk1.pcpi_mul_mul_2366_47_n_423 ,
       \genblk1.pcpi_mul_mul_2366_47_n_424 ,
       \genblk1.pcpi_mul_mul_2366_47_n_425 ,
       \genblk1.pcpi_mul_mul_2366_47_n_426 ,
       \genblk1.pcpi_mul_mul_2366_47_n_427 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_428 ,
       \genblk1.pcpi_mul_mul_2366_47_n_429 ,
       \genblk1.pcpi_mul_mul_2366_47_n_430 ,
       \genblk1.pcpi_mul_mul_2366_47_n_431 ,
       \genblk1.pcpi_mul_mul_2366_47_n_432 ,
       \genblk1.pcpi_mul_mul_2366_47_n_433 ,
       \genblk1.pcpi_mul_mul_2366_47_n_434 ,
       \genblk1.pcpi_mul_mul_2366_47_n_435 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_436 ,
       \genblk1.pcpi_mul_mul_2366_47_n_437 ,
       \genblk1.pcpi_mul_mul_2366_47_n_438 ,
       \genblk1.pcpi_mul_mul_2366_47_n_439 ,
       \genblk1.pcpi_mul_mul_2366_47_n_440 ,
       \genblk1.pcpi_mul_mul_2366_47_n_441 ,
       \genblk1.pcpi_mul_mul_2366_47_n_442 ,
       \genblk1.pcpi_mul_mul_2366_47_n_443 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_444 ,
       \genblk1.pcpi_mul_mul_2366_47_n_445 ,
       \genblk1.pcpi_mul_mul_2366_47_n_446 ,
       \genblk1.pcpi_mul_mul_2366_47_n_447 ,
       \genblk1.pcpi_mul_mul_2366_47_n_448 ,
       \genblk1.pcpi_mul_mul_2366_47_n_449 ,
       \genblk1.pcpi_mul_mul_2366_47_n_450 ,
       \genblk1.pcpi_mul_mul_2366_47_n_451 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_452 ,
       \genblk1.pcpi_mul_mul_2366_47_n_453 ,
       \genblk1.pcpi_mul_mul_2366_47_n_454 ,
       \genblk1.pcpi_mul_mul_2366_47_n_455 ,
       \genblk1.pcpi_mul_mul_2366_47_n_456 ,
       \genblk1.pcpi_mul_mul_2366_47_n_457 ,
       \genblk1.pcpi_mul_mul_2366_47_n_458 ,
       \genblk1.pcpi_mul_mul_2366_47_n_459 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_460 ,
       \genblk1.pcpi_mul_mul_2366_47_n_461 ,
       \genblk1.pcpi_mul_mul_2366_47_n_462 ,
       \genblk1.pcpi_mul_mul_2366_47_n_463 ,
       \genblk1.pcpi_mul_mul_2366_47_n_464 ,
       \genblk1.pcpi_mul_mul_2366_47_n_465 ,
       \genblk1.pcpi_mul_mul_2366_47_n_466 ,
       \genblk1.pcpi_mul_mul_2366_47_n_467 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_468 ,
       \genblk1.pcpi_mul_mul_2366_47_n_469 ,
       \genblk1.pcpi_mul_mul_2366_47_n_470 ,
       \genblk1.pcpi_mul_mul_2366_47_n_471 ,
       \genblk1.pcpi_mul_mul_2366_47_n_472 ,
       \genblk1.pcpi_mul_mul_2366_47_n_473 ,
       \genblk1.pcpi_mul_mul_2366_47_n_474 ,
       \genblk1.pcpi_mul_mul_2366_47_n_475 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_476 ,
       \genblk1.pcpi_mul_mul_2366_47_n_477 ,
       \genblk1.pcpi_mul_mul_2366_47_n_478 ,
       \genblk1.pcpi_mul_mul_2366_47_n_479 ,
       \genblk1.pcpi_mul_mul_2366_47_n_480 ,
       \genblk1.pcpi_mul_mul_2366_47_n_481 ,
       \genblk1.pcpi_mul_mul_2366_47_n_482 ,
       \genblk1.pcpi_mul_mul_2366_47_n_483 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_484 ,
       \genblk1.pcpi_mul_mul_2366_47_n_485 ,
       \genblk1.pcpi_mul_mul_2366_47_n_486 ,
       \genblk1.pcpi_mul_mul_2366_47_n_487 ,
       \genblk1.pcpi_mul_mul_2366_47_n_488 ,
       \genblk1.pcpi_mul_mul_2366_47_n_489 ,
       \genblk1.pcpi_mul_mul_2366_47_n_490 ,
       \genblk1.pcpi_mul_mul_2366_47_n_491 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_492 ,
       \genblk1.pcpi_mul_mul_2366_47_n_493 ,
       \genblk1.pcpi_mul_mul_2366_47_n_494 ,
       \genblk1.pcpi_mul_mul_2366_47_n_495 ,
       \genblk1.pcpi_mul_mul_2366_47_n_496 ,
       \genblk1.pcpi_mul_mul_2366_47_n_497 ,
       \genblk1.pcpi_mul_mul_2366_47_n_498 ,
       \genblk1.pcpi_mul_mul_2366_47_n_499 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_500 ,
       \genblk1.pcpi_mul_mul_2366_47_n_501 ,
       \genblk1.pcpi_mul_mul_2366_47_n_502 ,
       \genblk1.pcpi_mul_mul_2366_47_n_503 ,
       \genblk1.pcpi_mul_mul_2366_47_n_504 ,
       \genblk1.pcpi_mul_mul_2366_47_n_505 ,
       \genblk1.pcpi_mul_mul_2366_47_n_506 ,
       \genblk1.pcpi_mul_mul_2366_47_n_507 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_508 ,
       \genblk1.pcpi_mul_mul_2366_47_n_509 ,
       \genblk1.pcpi_mul_mul_2366_47_n_510 ,
       \genblk1.pcpi_mul_mul_2366_47_n_511 ,
       \genblk1.pcpi_mul_mul_2366_47_n_512 ,
       \genblk1.pcpi_mul_mul_2366_47_n_513 ,
       \genblk1.pcpi_mul_mul_2366_47_n_514 ,
       \genblk1.pcpi_mul_mul_2366_47_n_515 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_516 ,
       \genblk1.pcpi_mul_mul_2366_47_n_517 ,
       \genblk1.pcpi_mul_mul_2366_47_n_518 ,
       \genblk1.pcpi_mul_mul_2366_47_n_519 ,
       \genblk1.pcpi_mul_mul_2366_47_n_520 ,
       \genblk1.pcpi_mul_mul_2366_47_n_521 ,
       \genblk1.pcpi_mul_mul_2366_47_n_522 ,
       \genblk1.pcpi_mul_mul_2366_47_n_523 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_524 ,
       \genblk1.pcpi_mul_mul_2366_47_n_525 ,
       \genblk1.pcpi_mul_mul_2366_47_n_526 ,
       \genblk1.pcpi_mul_mul_2366_47_n_527 ,
       \genblk1.pcpi_mul_mul_2366_47_n_528 ,
       \genblk1.pcpi_mul_mul_2366_47_n_529 ,
       \genblk1.pcpi_mul_mul_2366_47_n_530 ,
       \genblk1.pcpi_mul_mul_2366_47_n_531 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_532 ,
       \genblk1.pcpi_mul_mul_2366_47_n_533 ,
       \genblk1.pcpi_mul_mul_2366_47_n_534 ,
       \genblk1.pcpi_mul_mul_2366_47_n_535 ,
       \genblk1.pcpi_mul_mul_2366_47_n_536 ,
       \genblk1.pcpi_mul_mul_2366_47_n_537 ,
       \genblk1.pcpi_mul_mul_2366_47_n_538 ,
       \genblk1.pcpi_mul_mul_2366_47_n_539 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_540 ,
       \genblk1.pcpi_mul_mul_2366_47_n_541 ,
       \genblk1.pcpi_mul_mul_2366_47_n_542 ,
       \genblk1.pcpi_mul_mul_2366_47_n_543 ,
       \genblk1.pcpi_mul_mul_2366_47_n_544 ,
       \genblk1.pcpi_mul_mul_2366_47_n_545 ,
       \genblk1.pcpi_mul_mul_2366_47_n_546 ,
       \genblk1.pcpi_mul_mul_2366_47_n_547 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_548 ,
       \genblk1.pcpi_mul_mul_2366_47_n_549 ,
       \genblk1.pcpi_mul_mul_2366_47_n_550 ,
       \genblk1.pcpi_mul_mul_2366_47_n_551 ,
       \genblk1.pcpi_mul_mul_2366_47_n_552 ,
       \genblk1.pcpi_mul_mul_2366_47_n_553 ,
       \genblk1.pcpi_mul_mul_2366_47_n_554 ,
       \genblk1.pcpi_mul_mul_2366_47_n_555 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_556 ,
       \genblk1.pcpi_mul_mul_2366_47_n_557 ,
       \genblk1.pcpi_mul_mul_2366_47_n_558 ,
       \genblk1.pcpi_mul_mul_2366_47_n_559 ,
       \genblk1.pcpi_mul_mul_2366_47_n_560 ,
       \genblk1.pcpi_mul_mul_2366_47_n_561 ,
       \genblk1.pcpi_mul_mul_2366_47_n_562 ,
       \genblk1.pcpi_mul_mul_2366_47_n_563 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_564 ,
       \genblk1.pcpi_mul_mul_2366_47_n_565 ,
       \genblk1.pcpi_mul_mul_2366_47_n_566 ,
       \genblk1.pcpi_mul_mul_2366_47_n_567 ,
       \genblk1.pcpi_mul_mul_2366_47_n_568 ,
       \genblk1.pcpi_mul_mul_2366_47_n_569 ,
       \genblk1.pcpi_mul_mul_2366_47_n_570 ,
       \genblk1.pcpi_mul_mul_2366_47_n_571 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_572 ,
       \genblk1.pcpi_mul_mul_2366_47_n_573 ,
       \genblk1.pcpi_mul_mul_2366_47_n_574 ,
       \genblk1.pcpi_mul_mul_2366_47_n_576 ,
       \genblk1.pcpi_mul_mul_2366_47_n_577 ,
       \genblk1.pcpi_mul_mul_2366_47_n_578 ,
       \genblk1.pcpi_mul_mul_2366_47_n_579 ,
       \genblk1.pcpi_mul_mul_2366_47_n_580 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_581 ,
       \genblk1.pcpi_mul_mul_2366_47_n_582 ,
       \genblk1.pcpi_mul_mul_2366_47_n_583 ,
       \genblk1.pcpi_mul_mul_2366_47_n_584 ,
       \genblk1.pcpi_mul_mul_2366_47_n_585 ,
       \genblk1.pcpi_mul_mul_2366_47_n_586 ,
       \genblk1.pcpi_mul_mul_2366_47_n_587 ,
       \genblk1.pcpi_mul_mul_2366_47_n_588 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_589 ,
       \genblk1.pcpi_mul_mul_2366_47_n_590 ,
       \genblk1.pcpi_mul_mul_2366_47_n_591 ,
       \genblk1.pcpi_mul_mul_2366_47_n_592 ,
       \genblk1.pcpi_mul_mul_2366_47_n_593 ,
       \genblk1.pcpi_mul_mul_2366_47_n_594 ,
       \genblk1.pcpi_mul_mul_2366_47_n_595 ,
       \genblk1.pcpi_mul_mul_2366_47_n_596 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_597 ,
       \genblk1.pcpi_mul_mul_2366_47_n_598 ,
       \genblk1.pcpi_mul_mul_2366_47_n_599 ,
       \genblk1.pcpi_mul_mul_2366_47_n_600 ,
       \genblk1.pcpi_mul_mul_2366_47_n_601 ,
       \genblk1.pcpi_mul_mul_2366_47_n_602 ,
       \genblk1.pcpi_mul_mul_2366_47_n_603 ,
       \genblk1.pcpi_mul_mul_2366_47_n_604 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_605 ,
       \genblk1.pcpi_mul_mul_2366_47_n_606 ,
       \genblk1.pcpi_mul_mul_2366_47_n_607 ,
       \genblk1.pcpi_mul_mul_2366_47_n_608 ,
       \genblk1.pcpi_mul_mul_2366_47_n_609 ,
       \genblk1.pcpi_mul_mul_2366_47_n_610 ,
       \genblk1.pcpi_mul_mul_2366_47_n_611 ,
       \genblk1.pcpi_mul_mul_2366_47_n_612 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_613 ,
       \genblk1.pcpi_mul_mul_2366_47_n_614 ,
       \genblk1.pcpi_mul_mul_2366_47_n_615 ,
       \genblk1.pcpi_mul_mul_2366_47_n_616 ,
       \genblk1.pcpi_mul_mul_2366_47_n_617 ,
       \genblk1.pcpi_mul_mul_2366_47_n_618 ,
       \genblk1.pcpi_mul_mul_2366_47_n_619 ,
       \genblk1.pcpi_mul_mul_2366_47_n_620 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_621 ,
       \genblk1.pcpi_mul_mul_2366_47_n_622 ,
       \genblk1.pcpi_mul_mul_2366_47_n_623 ,
       \genblk1.pcpi_mul_mul_2366_47_n_624 ,
       \genblk1.pcpi_mul_mul_2366_47_n_625 ,
       \genblk1.pcpi_mul_mul_2366_47_n_626 ,
       \genblk1.pcpi_mul_mul_2366_47_n_627 ,
       \genblk1.pcpi_mul_mul_2366_47_n_628 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_629 ,
       \genblk1.pcpi_mul_mul_2366_47_n_630 ,
       \genblk1.pcpi_mul_mul_2366_47_n_631 ,
       \genblk1.pcpi_mul_mul_2366_47_n_632 ,
       \genblk1.pcpi_mul_mul_2366_47_n_633 ,
       \genblk1.pcpi_mul_mul_2366_47_n_634 ,
       \genblk1.pcpi_mul_mul_2366_47_n_635 ,
       \genblk1.pcpi_mul_mul_2366_47_n_636 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_637 ,
       \genblk1.pcpi_mul_mul_2366_47_n_638 ,
       \genblk1.pcpi_mul_mul_2366_47_n_639 ,
       \genblk1.pcpi_mul_mul_2366_47_n_640 ,
       \genblk1.pcpi_mul_mul_2366_47_n_641 ,
       \genblk1.pcpi_mul_mul_2366_47_n_642 ,
       \genblk1.pcpi_mul_mul_2366_47_n_643 ,
       \genblk1.pcpi_mul_mul_2366_47_n_644 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_645 ,
       \genblk1.pcpi_mul_mul_2366_47_n_646 ,
       \genblk1.pcpi_mul_mul_2366_47_n_647 ,
       \genblk1.pcpi_mul_mul_2366_47_n_648 ,
       \genblk1.pcpi_mul_mul_2366_47_n_649 ,
       \genblk1.pcpi_mul_mul_2366_47_n_650 ,
       \genblk1.pcpi_mul_mul_2366_47_n_651 ,
       \genblk1.pcpi_mul_mul_2366_47_n_652 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_653 ,
       \genblk1.pcpi_mul_mul_2366_47_n_654 ,
       \genblk1.pcpi_mul_mul_2366_47_n_655 ,
       \genblk1.pcpi_mul_mul_2366_47_n_656 ,
       \genblk1.pcpi_mul_mul_2366_47_n_657 ,
       \genblk1.pcpi_mul_mul_2366_47_n_658 ,
       \genblk1.pcpi_mul_mul_2366_47_n_659 ,
       \genblk1.pcpi_mul_mul_2366_47_n_660 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_661 ,
       \genblk1.pcpi_mul_mul_2366_47_n_662 ,
       \genblk1.pcpi_mul_mul_2366_47_n_663 ,
       \genblk1.pcpi_mul_mul_2366_47_n_664 ,
       \genblk1.pcpi_mul_mul_2366_47_n_665 ,
       \genblk1.pcpi_mul_mul_2366_47_n_666 ,
       \genblk1.pcpi_mul_mul_2366_47_n_667 ,
       \genblk1.pcpi_mul_mul_2366_47_n_668 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_669 ,
       \genblk1.pcpi_mul_mul_2366_47_n_670 ,
       \genblk1.pcpi_mul_mul_2366_47_n_671 ,
       \genblk1.pcpi_mul_mul_2366_47_n_672 ,
       \genblk1.pcpi_mul_mul_2366_47_n_673 ,
       \genblk1.pcpi_mul_mul_2366_47_n_674 ,
       \genblk1.pcpi_mul_mul_2366_47_n_675 ,
       \genblk1.pcpi_mul_mul_2366_47_n_676 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_677 ,
       \genblk1.pcpi_mul_mul_2366_47_n_678 ,
       \genblk1.pcpi_mul_mul_2366_47_n_679 ,
       \genblk1.pcpi_mul_mul_2366_47_n_680 ,
       \genblk1.pcpi_mul_mul_2366_47_n_681 ,
       \genblk1.pcpi_mul_mul_2366_47_n_682 ,
       \genblk1.pcpi_mul_mul_2366_47_n_683 ,
       \genblk1.pcpi_mul_mul_2366_47_n_684 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_685 ,
       \genblk1.pcpi_mul_mul_2366_47_n_686 ,
       \genblk1.pcpi_mul_mul_2366_47_n_687 ,
       \genblk1.pcpi_mul_mul_2366_47_n_688 ,
       \genblk1.pcpi_mul_mul_2366_47_n_689 ,
       \genblk1.pcpi_mul_mul_2366_47_n_690 ,
       \genblk1.pcpi_mul_mul_2366_47_n_691 ,
       \genblk1.pcpi_mul_mul_2366_47_n_692 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_693 ,
       \genblk1.pcpi_mul_mul_2366_47_n_694 ,
       \genblk1.pcpi_mul_mul_2366_47_n_695 ,
       \genblk1.pcpi_mul_mul_2366_47_n_696 ,
       \genblk1.pcpi_mul_mul_2366_47_n_697 ,
       \genblk1.pcpi_mul_mul_2366_47_n_698 ,
       \genblk1.pcpi_mul_mul_2366_47_n_699 ,
       \genblk1.pcpi_mul_mul_2366_47_n_700 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_701 ,
       \genblk1.pcpi_mul_mul_2366_47_n_702 ,
       \genblk1.pcpi_mul_mul_2366_47_n_703 ,
       \genblk1.pcpi_mul_mul_2366_47_n_704 ,
       \genblk1.pcpi_mul_mul_2366_47_n_705 ,
       \genblk1.pcpi_mul_mul_2366_47_n_706 ,
       \genblk1.pcpi_mul_mul_2366_47_n_707 ,
       \genblk1.pcpi_mul_mul_2366_47_n_708 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_709 ,
       \genblk1.pcpi_mul_mul_2366_47_n_710 ,
       \genblk1.pcpi_mul_mul_2366_47_n_711 ,
       \genblk1.pcpi_mul_mul_2366_47_n_712 ,
       \genblk1.pcpi_mul_mul_2366_47_n_713 ,
       \genblk1.pcpi_mul_mul_2366_47_n_714 ,
       \genblk1.pcpi_mul_mul_2366_47_n_715 ,
       \genblk1.pcpi_mul_mul_2366_47_n_716 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_717 ,
       \genblk1.pcpi_mul_mul_2366_47_n_718 ,
       \genblk1.pcpi_mul_mul_2366_47_n_719 ,
       \genblk1.pcpi_mul_mul_2366_47_n_720 ,
       \genblk1.pcpi_mul_mul_2366_47_n_721 ,
       \genblk1.pcpi_mul_mul_2366_47_n_722 ,
       \genblk1.pcpi_mul_mul_2366_47_n_723 ,
       \genblk1.pcpi_mul_mul_2366_47_n_724 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_725 ,
       \genblk1.pcpi_mul_mul_2366_47_n_726 ,
       \genblk1.pcpi_mul_mul_2366_47_n_727 ,
       \genblk1.pcpi_mul_mul_2366_47_n_728 ,
       \genblk1.pcpi_mul_mul_2366_47_n_729 ,
       \genblk1.pcpi_mul_mul_2366_47_n_730 ,
       \genblk1.pcpi_mul_mul_2366_47_n_731 ,
       \genblk1.pcpi_mul_mul_2366_47_n_732 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_733 ,
       \genblk1.pcpi_mul_mul_2366_47_n_734 ,
       \genblk1.pcpi_mul_mul_2366_47_n_735 ,
       \genblk1.pcpi_mul_mul_2366_47_n_736 ,
       \genblk1.pcpi_mul_mul_2366_47_n_737 ,
       \genblk1.pcpi_mul_mul_2366_47_n_738 ,
       \genblk1.pcpi_mul_mul_2366_47_n_739 ,
       \genblk1.pcpi_mul_mul_2366_47_n_740 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_741 ,
       \genblk1.pcpi_mul_mul_2366_47_n_742 ,
       \genblk1.pcpi_mul_mul_2366_47_n_743 ,
       \genblk1.pcpi_mul_mul_2366_47_n_744 ,
       \genblk1.pcpi_mul_mul_2366_47_n_745 ,
       \genblk1.pcpi_mul_mul_2366_47_n_746 ,
       \genblk1.pcpi_mul_mul_2366_47_n_747 ,
       \genblk1.pcpi_mul_mul_2366_47_n_748 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_749 ,
       \genblk1.pcpi_mul_mul_2366_47_n_750 ,
       \genblk1.pcpi_mul_mul_2366_47_n_751 ,
       \genblk1.pcpi_mul_mul_2366_47_n_752 ,
       \genblk1.pcpi_mul_mul_2366_47_n_753 ,
       \genblk1.pcpi_mul_mul_2366_47_n_754 ,
       \genblk1.pcpi_mul_mul_2366_47_n_755 ,
       \genblk1.pcpi_mul_mul_2366_47_n_756 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_757 ,
       \genblk1.pcpi_mul_mul_2366_47_n_758 ,
       \genblk1.pcpi_mul_mul_2366_47_n_759 ,
       \genblk1.pcpi_mul_mul_2366_47_n_760 ,
       \genblk1.pcpi_mul_mul_2366_47_n_761 ,
       \genblk1.pcpi_mul_mul_2366_47_n_762 ,
       \genblk1.pcpi_mul_mul_2366_47_n_763 ,
       \genblk1.pcpi_mul_mul_2366_47_n_764 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_765 ,
       \genblk1.pcpi_mul_mul_2366_47_n_766 ,
       \genblk1.pcpi_mul_mul_2366_47_n_767 ,
       \genblk1.pcpi_mul_mul_2366_47_n_768 ,
       \genblk1.pcpi_mul_mul_2366_47_n_769 ,
       \genblk1.pcpi_mul_mul_2366_47_n_770 ,
       \genblk1.pcpi_mul_mul_2366_47_n_771 ,
       \genblk1.pcpi_mul_mul_2366_47_n_772 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_773 ,
       \genblk1.pcpi_mul_mul_2366_47_n_774 ,
       \genblk1.pcpi_mul_mul_2366_47_n_775 ,
       \genblk1.pcpi_mul_mul_2366_47_n_776 ,
       \genblk1.pcpi_mul_mul_2366_47_n_777 ,
       \genblk1.pcpi_mul_mul_2366_47_n_778 ,
       \genblk1.pcpi_mul_mul_2366_47_n_779 ,
       \genblk1.pcpi_mul_mul_2366_47_n_780 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_781 ,
       \genblk1.pcpi_mul_mul_2366_47_n_782 ,
       \genblk1.pcpi_mul_mul_2366_47_n_783 ,
       \genblk1.pcpi_mul_mul_2366_47_n_784 ,
       \genblk1.pcpi_mul_mul_2366_47_n_785 ,
       \genblk1.pcpi_mul_mul_2366_47_n_786 ,
       \genblk1.pcpi_mul_mul_2366_47_n_787 ,
       \genblk1.pcpi_mul_mul_2366_47_n_788 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_789 ,
       \genblk1.pcpi_mul_mul_2366_47_n_790 ,
       \genblk1.pcpi_mul_mul_2366_47_n_791 ,
       \genblk1.pcpi_mul_mul_2366_47_n_792 ,
       \genblk1.pcpi_mul_mul_2366_47_n_793 ,
       \genblk1.pcpi_mul_mul_2366_47_n_794 ,
       \genblk1.pcpi_mul_mul_2366_47_n_795 ,
       \genblk1.pcpi_mul_mul_2366_47_n_796 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_797 ,
       \genblk1.pcpi_mul_mul_2366_47_n_798 ,
       \genblk1.pcpi_mul_mul_2366_47_n_799 ,
       \genblk1.pcpi_mul_mul_2366_47_n_800 ,
       \genblk1.pcpi_mul_mul_2366_47_n_801 ,
       \genblk1.pcpi_mul_mul_2366_47_n_802 ,
       \genblk1.pcpi_mul_mul_2366_47_n_803 ,
       \genblk1.pcpi_mul_mul_2366_47_n_804 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_805 ,
       \genblk1.pcpi_mul_mul_2366_47_n_806 ,
       \genblk1.pcpi_mul_mul_2366_47_n_807 ,
       \genblk1.pcpi_mul_mul_2366_47_n_808 ,
       \genblk1.pcpi_mul_mul_2366_47_n_809 ,
       \genblk1.pcpi_mul_mul_2366_47_n_810 ,
       \genblk1.pcpi_mul_mul_2366_47_n_811 ,
       \genblk1.pcpi_mul_mul_2366_47_n_812 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_813 ,
       \genblk1.pcpi_mul_mul_2366_47_n_814 ,
       \genblk1.pcpi_mul_mul_2366_47_n_815 ,
       \genblk1.pcpi_mul_mul_2366_47_n_816 ,
       \genblk1.pcpi_mul_mul_2366_47_n_817 ,
       \genblk1.pcpi_mul_mul_2366_47_n_818 ,
       \genblk1.pcpi_mul_mul_2366_47_n_819 ,
       \genblk1.pcpi_mul_mul_2366_47_n_820 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_821 ,
       \genblk1.pcpi_mul_mul_2366_47_n_822 ,
       \genblk1.pcpi_mul_mul_2366_47_n_823 ,
       \genblk1.pcpi_mul_mul_2366_47_n_824 ,
       \genblk1.pcpi_mul_mul_2366_47_n_825 ,
       \genblk1.pcpi_mul_mul_2366_47_n_826 ,
       \genblk1.pcpi_mul_mul_2366_47_n_827 ,
       \genblk1.pcpi_mul_mul_2366_47_n_828 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_829 ,
       \genblk1.pcpi_mul_mul_2366_47_n_830 ,
       \genblk1.pcpi_mul_mul_2366_47_n_831 ,
       \genblk1.pcpi_mul_mul_2366_47_n_832 ,
       \genblk1.pcpi_mul_mul_2366_47_n_833 ,
       \genblk1.pcpi_mul_mul_2366_47_n_834 ,
       \genblk1.pcpi_mul_mul_2366_47_n_835 ,
       \genblk1.pcpi_mul_mul_2366_47_n_836 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_837 ,
       \genblk1.pcpi_mul_mul_2366_47_n_838 ,
       \genblk1.pcpi_mul_mul_2366_47_n_839 ,
       \genblk1.pcpi_mul_mul_2366_47_n_840 ,
       \genblk1.pcpi_mul_mul_2366_47_n_841 ,
       \genblk1.pcpi_mul_mul_2366_47_n_842 ,
       \genblk1.pcpi_mul_mul_2366_47_n_843 ,
       \genblk1.pcpi_mul_mul_2366_47_n_844 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_845 ,
       \genblk1.pcpi_mul_mul_2366_47_n_846 ,
       \genblk1.pcpi_mul_mul_2366_47_n_847 ,
       \genblk1.pcpi_mul_mul_2366_47_n_848 ,
       \genblk1.pcpi_mul_mul_2366_47_n_849 ,
       \genblk1.pcpi_mul_mul_2366_47_n_850 ,
       \genblk1.pcpi_mul_mul_2366_47_n_851 ,
       \genblk1.pcpi_mul_mul_2366_47_n_852 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_853 ,
       \genblk1.pcpi_mul_mul_2366_47_n_854 ,
       \genblk1.pcpi_mul_mul_2366_47_n_855 ,
       \genblk1.pcpi_mul_mul_2366_47_n_856 ,
       \genblk1.pcpi_mul_mul_2366_47_n_857 ,
       \genblk1.pcpi_mul_mul_2366_47_n_858 ,
       \genblk1.pcpi_mul_mul_2366_47_n_859 ,
       \genblk1.pcpi_mul_mul_2366_47_n_860 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_861 ,
       \genblk1.pcpi_mul_mul_2366_47_n_862 ,
       \genblk1.pcpi_mul_mul_2366_47_n_863 ,
       \genblk1.pcpi_mul_mul_2366_47_n_864 ,
       \genblk1.pcpi_mul_mul_2366_47_n_865 ,
       \genblk1.pcpi_mul_mul_2366_47_n_866 ,
       \genblk1.pcpi_mul_mul_2366_47_n_867 ,
       \genblk1.pcpi_mul_mul_2366_47_n_868 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_869 ,
       \genblk1.pcpi_mul_mul_2366_47_n_870 ,
       \genblk1.pcpi_mul_mul_2366_47_n_871 ,
       \genblk1.pcpi_mul_mul_2366_47_n_872 ,
       \genblk1.pcpi_mul_mul_2366_47_n_873 ,
       \genblk1.pcpi_mul_mul_2366_47_n_874 ,
       \genblk1.pcpi_mul_mul_2366_47_n_875 ,
       \genblk1.pcpi_mul_mul_2366_47_n_876 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_877 ,
       \genblk1.pcpi_mul_mul_2366_47_n_878 ,
       \genblk1.pcpi_mul_mul_2366_47_n_879 ,
       \genblk1.pcpi_mul_mul_2366_47_n_880 ,
       \genblk1.pcpi_mul_mul_2366_47_n_881 ,
       \genblk1.pcpi_mul_mul_2366_47_n_882 ,
       \genblk1.pcpi_mul_mul_2366_47_n_883 ,
       \genblk1.pcpi_mul_mul_2366_47_n_884 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_885 ,
       \genblk1.pcpi_mul_mul_2366_47_n_886 ,
       \genblk1.pcpi_mul_mul_2366_47_n_887 ,
       \genblk1.pcpi_mul_mul_2366_47_n_888 ,
       \genblk1.pcpi_mul_mul_2366_47_n_889 ,
       \genblk1.pcpi_mul_mul_2366_47_n_890 ,
       \genblk1.pcpi_mul_mul_2366_47_n_891 ,
       \genblk1.pcpi_mul_mul_2366_47_n_892 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_893 ,
       \genblk1.pcpi_mul_mul_2366_47_n_894 ,
       \genblk1.pcpi_mul_mul_2366_47_n_895 ,
       \genblk1.pcpi_mul_mul_2366_47_n_896 ,
       \genblk1.pcpi_mul_mul_2366_47_n_897 ,
       \genblk1.pcpi_mul_mul_2366_47_n_898 ,
       \genblk1.pcpi_mul_mul_2366_47_n_899 ,
       \genblk1.pcpi_mul_mul_2366_47_n_900 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_901 ,
       \genblk1.pcpi_mul_mul_2366_47_n_902 ,
       \genblk1.pcpi_mul_mul_2366_47_n_903 ,
       \genblk1.pcpi_mul_mul_2366_47_n_904 ,
       \genblk1.pcpi_mul_mul_2366_47_n_905 ,
       \genblk1.pcpi_mul_mul_2366_47_n_906 ,
       \genblk1.pcpi_mul_mul_2366_47_n_907 ,
       \genblk1.pcpi_mul_mul_2366_47_n_908 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_909 ,
       \genblk1.pcpi_mul_mul_2366_47_n_910 ,
       \genblk1.pcpi_mul_mul_2366_47_n_911 ,
       \genblk1.pcpi_mul_mul_2366_47_n_912 ,
       \genblk1.pcpi_mul_mul_2366_47_n_913 ,
       \genblk1.pcpi_mul_mul_2366_47_n_914 ,
       \genblk1.pcpi_mul_mul_2366_47_n_915 ,
       \genblk1.pcpi_mul_mul_2366_47_n_916 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_917 ,
       \genblk1.pcpi_mul_mul_2366_47_n_918 ,
       \genblk1.pcpi_mul_mul_2366_47_n_919 ,
       \genblk1.pcpi_mul_mul_2366_47_n_920 ,
       \genblk1.pcpi_mul_mul_2366_47_n_921 ,
       \genblk1.pcpi_mul_mul_2366_47_n_922 ,
       \genblk1.pcpi_mul_mul_2366_47_n_923 ,
       \genblk1.pcpi_mul_mul_2366_47_n_924 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_925 ,
       \genblk1.pcpi_mul_mul_2366_47_n_926 ,
       \genblk1.pcpi_mul_mul_2366_47_n_927 ,
       \genblk1.pcpi_mul_mul_2366_47_n_928 ,
       \genblk1.pcpi_mul_mul_2366_47_n_929 ,
       \genblk1.pcpi_mul_mul_2366_47_n_930 ,
       \genblk1.pcpi_mul_mul_2366_47_n_931 ,
       \genblk1.pcpi_mul_mul_2366_47_n_932 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_933 ,
       \genblk1.pcpi_mul_mul_2366_47_n_934 ,
       \genblk1.pcpi_mul_mul_2366_47_n_935 ,
       \genblk1.pcpi_mul_mul_2366_47_n_936 ,
       \genblk1.pcpi_mul_mul_2366_47_n_937 ,
       \genblk1.pcpi_mul_mul_2366_47_n_938 ,
       \genblk1.pcpi_mul_mul_2366_47_n_939 ,
       \genblk1.pcpi_mul_mul_2366_47_n_940 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_941 ,
       \genblk1.pcpi_mul_mul_2366_47_n_942 ,
       \genblk1.pcpi_mul_mul_2366_47_n_943 ,
       \genblk1.pcpi_mul_mul_2366_47_n_944 ,
       \genblk1.pcpi_mul_mul_2366_47_n_945 ,
       \genblk1.pcpi_mul_mul_2366_47_n_946 ,
       \genblk1.pcpi_mul_mul_2366_47_n_947 ,
       \genblk1.pcpi_mul_mul_2366_47_n_948 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_949 ,
       \genblk1.pcpi_mul_mul_2366_47_n_950 ,
       \genblk1.pcpi_mul_mul_2366_47_n_951 ,
       \genblk1.pcpi_mul_mul_2366_47_n_952 ,
       \genblk1.pcpi_mul_mul_2366_47_n_953 ,
       \genblk1.pcpi_mul_mul_2366_47_n_954 ,
       \genblk1.pcpi_mul_mul_2366_47_n_955 ,
       \genblk1.pcpi_mul_mul_2366_47_n_956 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_957 ,
       \genblk1.pcpi_mul_mul_2366_47_n_958 ,
       \genblk1.pcpi_mul_mul_2366_47_n_959 ,
       \genblk1.pcpi_mul_mul_2366_47_n_960 ,
       \genblk1.pcpi_mul_mul_2366_47_n_961 ,
       \genblk1.pcpi_mul_mul_2366_47_n_962 ,
       \genblk1.pcpi_mul_mul_2366_47_n_963 ,
       \genblk1.pcpi_mul_mul_2366_47_n_964 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_965 ,
       \genblk1.pcpi_mul_mul_2366_47_n_966 ,
       \genblk1.pcpi_mul_mul_2366_47_n_967 ,
       \genblk1.pcpi_mul_mul_2366_47_n_968 ,
       \genblk1.pcpi_mul_mul_2366_47_n_969 ,
       \genblk1.pcpi_mul_mul_2366_47_n_970 ,
       \genblk1.pcpi_mul_mul_2366_47_n_971 ,
       \genblk1.pcpi_mul_mul_2366_47_n_972 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_973 ,
       \genblk1.pcpi_mul_mul_2366_47_n_974 ,
       \genblk1.pcpi_mul_mul_2366_47_n_975 ,
       \genblk1.pcpi_mul_mul_2366_47_n_976 ,
       \genblk1.pcpi_mul_mul_2366_47_n_977 ,
       \genblk1.pcpi_mul_mul_2366_47_n_978 ,
       \genblk1.pcpi_mul_mul_2366_47_n_979 ,
       \genblk1.pcpi_mul_mul_2366_47_n_980 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_981 ,
       \genblk1.pcpi_mul_mul_2366_47_n_982 ,
       \genblk1.pcpi_mul_mul_2366_47_n_983 ,
       \genblk1.pcpi_mul_mul_2366_47_n_984 ,
       \genblk1.pcpi_mul_mul_2366_47_n_985 ,
       \genblk1.pcpi_mul_mul_2366_47_n_986 ,
       \genblk1.pcpi_mul_mul_2366_47_n_987 ,
       \genblk1.pcpi_mul_mul_2366_47_n_988 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_989 ,
       \genblk1.pcpi_mul_mul_2366_47_n_990 ,
       \genblk1.pcpi_mul_mul_2366_47_n_991 ,
       \genblk1.pcpi_mul_mul_2366_47_n_992 ,
       \genblk1.pcpi_mul_mul_2366_47_n_993 ,
       \genblk1.pcpi_mul_mul_2366_47_n_994 ,
       \genblk1.pcpi_mul_mul_2366_47_n_995 ,
       \genblk1.pcpi_mul_mul_2366_47_n_996 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_997 ,
       \genblk1.pcpi_mul_mul_2366_47_n_998 ,
       \genblk1.pcpi_mul_mul_2366_47_n_999 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1000 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1001 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1002 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1003 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1004 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1005 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1006 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1007 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1008 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1009 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1010 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1011 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1012 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1013 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1014 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1015 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1016 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1017 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1018 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1019 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1020 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1021 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1022 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1023 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1024 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1025 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1026 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1027 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1028 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1029 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1030 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1031 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1032 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1033 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1034 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1035 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1036 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1037 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1038 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1039 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1040 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1041 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1042 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1043 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1044 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1045 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1046 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1047 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1048 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1049 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1050 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1051 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1052 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1053 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1054 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1055 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1056 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1057 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1058 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1059 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1060 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1061 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1062 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1063 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1064 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1065 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1066 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1067 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1068 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1069 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1070 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1071 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1072 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1073 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1074 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1075 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1076 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1077 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1078 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1079 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1080 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1081 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1082 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1083 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1084 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1085 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1086 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1087 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1088 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1089 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1090 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1091 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1092 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1093 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1094 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1095 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1096 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1097 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1098 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1099 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1100 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1101 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1102 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1103 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1104 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1105 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1106 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1107 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1108 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1109 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1110 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1111 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1112 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1113 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1114 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1115 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1116 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1117 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1118 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1119 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1120 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1121 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1122 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1123 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1124 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1125 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1126 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1127 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1128 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1129 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1130 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1131 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1132 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1133 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1134 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1135 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1136 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1137 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1138 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1139 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1140 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1141 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1142 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1143 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1144 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1145 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1146 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1147 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1148 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1149 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1150 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1151 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1152 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1153 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1154 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1155 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1156 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1157 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1158 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1159 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1160 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1161 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1162 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1163 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1164 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1165 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1166 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1167 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1168 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1169 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1170 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1171 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1172 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1173 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1174 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1175 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1176 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1177 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1178 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1179 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1180 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1181 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1182 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1183 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1184 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1185 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1186 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1187 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1188 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1189 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1190 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1191 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1192 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1193 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1194 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1195 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1196 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1197 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1198 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1199 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1200 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1201 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1202 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1203 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1204 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1205 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1206 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1207 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1208 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1209 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1210 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1211 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1212 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1213 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1214 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1215 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1216 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1217 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1218 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1219 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1220 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1221 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1222 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1223 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1224 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1225 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1226 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1227 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1228 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1229 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1230 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1231 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1232 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1233 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1234 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1235 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1236 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1237 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1238 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1239 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1240 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1241 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1242 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1243 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1244 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1245 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1246 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1247 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1248 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1249 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1250 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1251 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1252 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1253 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1254 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1255 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1256 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1257 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1258 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1259 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1260 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1261 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1262 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1263 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1264 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1265 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1266 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1267 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1268 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1269 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1270 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1271 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1272 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1273 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1274 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1275 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1276 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1277 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1278 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1279 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1280 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1281 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1282 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1283 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1284 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1285 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1286 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1287 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1288 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1289 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1290 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1291 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1292 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1293 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1294 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1295 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1296 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1297 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1298 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1299 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1300 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1301 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1302 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1303 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1304 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1305 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1306 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1307 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1308 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1309 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1310 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1311 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1312 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1313 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1314 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1315 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1316 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1317 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1318 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1319 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1320 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1321 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1322 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1323 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1324 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1325 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1326 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1327 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1328 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1329 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1330 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1331 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1332 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1333 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1334 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1335 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1336 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1337 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1338 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1339 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1340 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1341 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1342 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1343 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1344 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1345 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1346 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1347 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1348 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1349 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1350 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1351 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1352 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1353 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1354 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1355 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1356 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1357 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1358 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1359 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1360 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1361 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1362 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1363 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1364 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1365 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1366 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1367 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1368 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1369 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1370 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1371 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1372 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1373 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1374 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1375 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1376 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1377 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1378 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1379 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1380 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1381 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1382 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1383 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1384 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1385 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1386 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1387 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1388 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1389 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1390 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1391 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1392 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1393 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1394 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1395 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1396 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1397 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1398 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1399 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1400 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1401 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1402 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1403 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1404 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1405 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1406 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1407 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1408 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1409 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1410 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1411 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1412 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1413 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1414 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1415 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1416 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1417 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1418 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1419 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1420 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1421 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1422 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1423 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1424 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1425 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1426 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1427 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1428 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1429 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1430 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1431 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1432 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1433 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1434 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1435 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1436 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1437 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1438 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1439 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1440 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1441 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1442 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1443 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1444 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1445 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1446 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1447 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1448 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1449 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1450 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1451 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1453 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1454 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1455 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1456 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1457 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1458 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1459 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1460 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1461 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1462 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1463 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1464 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1465 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1466 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1467 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1468 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1469 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1470 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1471 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1472 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1473 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1474 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1475 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1476 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1477 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1478 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1479 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1480 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1481 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1482 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1483 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1484 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1485 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1486 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1487 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1488 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1489 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1490 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1491 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1492 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1493 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1494 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1495 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1496 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1497 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1498 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1499 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1500 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1501 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1502 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1503 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1504 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1505 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1506 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1507 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1508 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1509 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1510 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1511 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1512 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1513 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1514 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1515 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1516 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1517 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1518 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1519 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1520 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1521 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1522 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1523 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1524 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1525 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1526 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1527 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1528 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1529 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1530 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1531 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1532 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1533 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1534 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1535 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1536 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1537 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1538 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1539 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1540 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1541 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1542 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1543 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1544 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1545 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1546 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1547 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1548 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1549 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1550 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1551 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1552 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1553 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1554 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1555 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1556 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1557 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1558 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1559 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1560 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1561 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1562 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1563 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1564 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1565 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1566 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1567 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1568 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1569 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1570 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1571 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1572 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1573 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1574 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1575 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1576 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1577 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1578 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1579 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1580 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1581 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1582 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1583 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1584 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1585 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1586 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1587 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1588 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1589 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1590 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1591 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1592 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1593 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1594 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1595 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1596 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1597 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1598 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1599 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1600 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1601 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1602 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1603 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1604 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1605 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1606 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1607 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1608 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1609 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1610 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1611 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1612 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1613 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1614 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1615 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1616 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1617 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1618 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1619 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1620 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1621 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1622 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1623 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1624 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1625 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1626 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1627 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1628 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1629 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1631 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1632 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1633 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1634 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1635 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1636 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1637 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1638 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1639 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1640 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1641 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1642 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1643 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1644 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1645 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1646 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1647 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1648 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1649 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1650 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1651 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1652 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1653 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1654 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1655 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1656 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1657 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1658 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1659 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1660 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1661 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1662 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1663 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1664 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1665 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1666 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1667 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1668 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1669 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1670 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1671 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1672 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1673 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1674 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1675 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1676 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1677 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1678 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1679 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1680 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1681 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1682 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1683 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1684 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1685 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1686 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1687 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1688 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1689 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1690 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1691 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1692 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1693 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1694 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1695 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1696 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1697 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1698 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1699 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1700 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1701 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1702 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1703 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1704 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1705 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1706 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1707 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1708 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1709 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1710 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1711 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1712 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1713 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1714 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1715 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1716 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1717 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1718 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1719 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1720 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1721 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1722 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1723 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1724 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1725 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1726 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1727 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1728 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1729 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1730 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1731 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1732 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1733 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1734 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1735 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1736 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1737 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1738 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1739 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1740 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1741 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1742 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1743 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1744 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1745 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1746 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1747 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1748 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1749 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1750 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1751 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1752 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1753 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1754 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1755 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1756 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1757 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1758 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1759 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1760 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1761 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1762 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1763 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1764 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1765 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1766 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1767 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1768 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1769 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1770 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1771 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1772 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1773 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1774 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1775 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1776 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1777 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1778 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1779 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1780 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1781 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1782 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1783 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1784 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1785 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1786 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1787 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1788 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1789 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1790 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1791 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1792 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1793 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1794 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1795 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1796 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1797 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1798 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1799 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1800 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1801 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1802 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1803 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1804 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1805 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1806 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1807 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1808 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1809 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1810 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1811 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1812 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1813 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1814 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1815 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1816 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1817 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1818 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1819 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1820 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1821 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1822 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1823 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1824 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1825 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1827 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1828 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1829 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1830 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1831 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1832 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1833 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1834 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1835 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1836 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1837 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1838 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1839 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1840 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1841 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1842 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1843 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1844 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1845 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1846 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1847 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1848 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1849 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1850 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1851 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1852 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1853 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1854 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1855 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1856 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1857 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1858 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1859 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1860 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1861 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1862 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1863 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1864 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1865 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1866 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1867 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1868 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1869 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1870 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1871 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1872 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1873 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1874 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1875 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1876 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1877 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1878 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1879 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1880 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1881 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1882 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1883 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1884 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1885 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1886 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1887 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1888 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1889 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1890 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1891 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1892 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1893 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1894 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1895 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1896 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1897 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1898 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1899 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1900 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1901 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1902 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1903 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1904 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1905 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1906 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1907 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1908 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1909 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1910 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1911 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1912 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1913 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1914 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1915 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1916 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1917 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1918 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1920 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1921 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1922 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1923 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1924 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1925 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1926 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1927 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1928 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1929 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1930 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1931 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1932 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1933 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1934 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1935 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1936 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1937 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1938 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1939 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1940 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1941 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1942 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1943 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1944 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1945 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1946 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1947 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1948 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1949 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1950 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1951 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1952 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1953 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1954 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1955 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1956 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1957 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1958 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1959 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1960 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1961 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1962 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1963 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1964 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1965 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1966 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1967 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1968 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1969 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1970 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1971 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1972 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1973 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1974 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1975 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1976 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1977 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1978 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1979 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1980 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1981 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1982 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1983 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1984 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1985 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1986 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1987 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1988 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1989 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1990 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1991 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1992 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_1993 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1994 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1995 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1996 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1997 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1998 ,
       \genblk1.pcpi_mul_mul_2366_47_n_1999 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2000 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2001 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2002 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2003 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2004 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2005 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2006 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2007 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2008 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2009 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2010 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2011 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2012 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2013 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2014 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2015 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2016 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2017 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2018 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2019 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2020 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2021 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2022 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2023 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2024 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2025 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2026 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2027 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2028 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2029 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2030 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2031 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2032 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2033 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2034 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2035 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2036 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2037 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2038 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2039 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2040 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2041 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2042 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2043 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2044 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2045 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2046 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2047 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2048 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2049 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2050 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2051 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2052 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2053 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2054 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2055 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2056 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2057 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2058 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2059 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2060 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2061 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2062 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2063 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2064 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2065 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2066 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2067 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2068 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2069 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2070 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2071 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2072 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2073 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2074 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2075 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2076 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2077 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2078 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2079 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2080 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2081 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2082 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2083 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2084 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2085 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2086 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2087 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2088 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2090 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2091 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2092 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2093 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2094 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2095 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2096 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2097 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2098 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2099 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2100 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2101 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2102 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2103 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2104 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2105 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2106 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2107 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2108 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2109 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2110 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2111 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2112 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2113 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2114 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2115 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2116 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2117 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2118 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2119 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2120 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2121 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2122 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2123 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2124 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2125 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2126 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2127 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2128 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2129 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2130 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2131 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2132 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2133 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2134 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2135 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2136 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2137 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2138 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2139 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2140 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2141 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2142 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2143 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2144 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2145 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2146 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2147 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2148 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2149 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2150 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2151 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2152 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2153 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2154 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2155 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2156 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2157 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2158 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2159 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2160 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2161 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2162 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2163 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2164 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2165 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2166 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2167 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2168 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2169 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2170 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2171 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2172 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2173 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2174 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2175 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2176 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2177 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2178 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2179 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2180 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2181 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2182 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2183 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2184 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2185 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2186 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2187 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2188 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2190 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2191 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2192 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2193 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2194 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2195 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2196 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2197 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2198 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2199 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2200 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2201 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2202 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2203 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2204 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2205 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2206 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2207 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2208 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2209 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2210 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2211 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2212 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2213 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2214 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2215 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2216 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2217 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2218 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2219 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2220 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2221 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2222 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2223 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2224 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2225 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2226 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2227 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2228 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2229 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2230 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2231 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2232 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2233 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2234 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2235 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2236 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2237 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2238 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2239 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2240 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2241 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2242 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2243 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2244 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2245 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2246 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2247 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2248 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2249 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2250 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2251 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2252 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2253 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2254 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2255 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2256 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2257 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2258 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2259 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2260 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2261 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2262 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2263 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2264 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2265 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2266 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2267 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2268 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2269 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2270 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2272 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2273 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2274 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2275 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2276 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2277 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2278 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2279 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2280 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2281 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2282 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2283 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2284 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2285 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2286 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2287 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2288 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2289 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2290 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2291 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2292 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2293 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2294 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2295 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2296 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2297 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2298 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2299 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2300 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2301 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2302 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2303 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2304 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2305 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2306 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2307 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2308 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2309 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2310 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2311 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2312 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2313 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2314 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2315 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2316 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2317 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2318 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2319 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2320 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2321 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2322 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2323 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2324 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2325 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2326 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2327 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2328 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2329 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2330 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2332 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2333 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2334 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2335 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2336 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2337 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2338 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2339 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2340 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2341 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2342 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2343 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2344 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2345 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2346 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2347 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2348 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2349 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2350 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2351 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2352 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2353 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2354 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2355 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2356 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2357 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2358 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2359 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2360 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2361 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2362 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2363 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2364 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2365 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2366 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2367 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2368 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2369 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2370 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2371 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2372 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2373 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2374 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2375 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2376 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2377 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2378 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2379 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2380 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2382 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2383 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2384 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2385 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2386 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2387 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2388 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2389 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2390 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2391 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2392 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2393 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2394 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2395 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2396 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2397 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2398 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2399 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2400 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2401 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2402 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2403 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2404 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2405 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2406 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2407 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2408 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2410 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2411 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2412 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2413 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2414 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2415 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2416 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2417 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2418 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2419 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2420 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2421 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2422 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2423 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2424 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2425 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2426 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2427 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2428 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2429 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2430 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2431 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2432 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2433 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2434 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2435 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2436 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2438 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2439 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2440 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2441 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2442 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2444 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2446 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2448 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2450 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2452 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2454 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2456 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2458 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2460 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2462 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2464 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2466 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2468 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2470 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2472 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2474 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2476 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2478 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2480 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2482 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2484 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2486 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2488 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2490 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2492 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2494 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2496 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2498 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2500 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2502 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2504 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2506 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2508 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2510 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2512 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2514 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2516 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2518 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2520 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2522 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2524 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2526 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2528 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2530 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2532 ;
  wire \genblk1.pcpi_mul_mul_2366_47_n_2534 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2536 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2538 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2540 ,
       \genblk1.pcpi_mul_mul_2366_47_n_2542 , \genblk1.pcpi_mul_n_91 ,
       \genblk1.pcpi_mul_n_92 , \genblk1.pcpi_mul_n_93 ;
  wire \genblk1.pcpi_mul_n_94 , \genblk1.pcpi_mul_n_95 ,
       \genblk1.pcpi_mul_n_96 , \genblk1.pcpi_mul_n_97 ,
       \genblk1.pcpi_mul_n_98 , \genblk1.pcpi_mul_n_99 ,
       \genblk1.pcpi_mul_n_100 , \genblk1.pcpi_mul_n_101 ;
  wire \genblk1.pcpi_mul_n_102 , \genblk1.pcpi_mul_n_103 ,
       \genblk1.pcpi_mul_n_104 , \genblk1.pcpi_mul_n_105 ,
       \genblk1.pcpi_mul_n_106 , \genblk1.pcpi_mul_n_107 ,
       \genblk1.pcpi_mul_n_108 , \genblk1.pcpi_mul_n_109 ;
  wire \genblk1.pcpi_mul_n_110 , \genblk1.pcpi_mul_n_111 ,
       \genblk1.pcpi_mul_n_112 , \genblk1.pcpi_mul_n_113 ,
       \genblk1.pcpi_mul_n_114 , \genblk1.pcpi_mul_n_115 ,
       \genblk1.pcpi_mul_n_116 , \genblk1.pcpi_mul_n_117 ;
  wire \genblk1.pcpi_mul_n_118 , \genblk1.pcpi_mul_n_119 ,
       \genblk1.pcpi_mul_n_120 , \genblk1.pcpi_mul_n_121 ,
       \genblk1.pcpi_mul_n_122 , \genblk1.pcpi_mul_n_123 ,
       \genblk1.pcpi_mul_n_124 , \genblk1.pcpi_mul_n_125 ;
  wire \genblk1.pcpi_mul_n_126 , \genblk1.pcpi_mul_n_127 ,
       \genblk1.pcpi_mul_n_128 , \genblk1.pcpi_mul_n_129 ,
       \genblk1.pcpi_mul_n_130 , \genblk1.pcpi_mul_n_131 ,
       \genblk1.pcpi_mul_n_132 , \genblk1.pcpi_mul_n_133 ;
  wire \genblk1.pcpi_mul_n_134 , \genblk1.pcpi_mul_n_135 ,
       \genblk1.pcpi_mul_n_136 , \genblk1.pcpi_mul_n_137 ,
       \genblk1.pcpi_mul_n_138 , \genblk1.pcpi_mul_n_139 ,
       \genblk1.pcpi_mul_n_140 , \genblk1.pcpi_mul_n_141 ;
  wire \genblk1.pcpi_mul_n_142 , \genblk1.pcpi_mul_n_143 ,
       \genblk1.pcpi_mul_n_144 , \genblk1.pcpi_mul_n_145 ,
       \genblk1.pcpi_mul_n_146 , \genblk1.pcpi_mul_n_147 ,
       \genblk1.pcpi_mul_n_148 , \genblk1.pcpi_mul_n_149 ;
  wire \genblk1.pcpi_mul_n_150 , \genblk1.pcpi_mul_n_151 ,
       \genblk1.pcpi_mul_n_152 , \genblk1.pcpi_mul_n_153 ,
       \genblk1.pcpi_mul_n_154 , \genblk1.pcpi_mul_shift_out ,
       \genblk2.pcpi_div_instr_div , \genblk2.pcpi_div_instr_divu ;
  wire \genblk2.pcpi_div_instr_rem , \genblk2.pcpi_div_instr_remu ,
       \genblk2.pcpi_div_lte_2493_16_n_0 ,
       \genblk2.pcpi_div_lte_2493_16_n_1 ,
       \genblk2.pcpi_div_lte_2493_16_n_2 ,
       \genblk2.pcpi_div_lte_2493_16_n_3 ,
       \genblk2.pcpi_div_lte_2493_16_n_4 ,
       \genblk2.pcpi_div_lte_2493_16_n_5 ;
  wire \genblk2.pcpi_div_lte_2493_16_n_6 ,
       \genblk2.pcpi_div_lte_2493_16_n_7 ,
       \genblk2.pcpi_div_lte_2493_16_n_8 ,
       \genblk2.pcpi_div_lte_2493_16_n_9 ,
       \genblk2.pcpi_div_lte_2493_16_n_10 ,
       \genblk2.pcpi_div_lte_2493_16_n_11 ,
       \genblk2.pcpi_div_lte_2493_16_n_12 ,
       \genblk2.pcpi_div_lte_2493_16_n_13 ;
  wire \genblk2.pcpi_div_lte_2493_16_n_14 ,
       \genblk2.pcpi_div_lte_2493_16_n_15 ,
       \genblk2.pcpi_div_lte_2493_16_n_16 ,
       \genblk2.pcpi_div_lte_2493_16_n_17 ,
       \genblk2.pcpi_div_lte_2493_16_n_18 ,
       \genblk2.pcpi_div_lte_2493_16_n_19 ,
       \genblk2.pcpi_div_lte_2493_16_n_20 ,
       \genblk2.pcpi_div_lte_2493_16_n_21 ;
  wire \genblk2.pcpi_div_lte_2493_16_n_22 ,
       \genblk2.pcpi_div_lte_2493_16_n_23 ,
       \genblk2.pcpi_div_lte_2493_16_n_24 ,
       \genblk2.pcpi_div_lte_2493_16_n_25 ,
       \genblk2.pcpi_div_lte_2493_16_n_26 ,
       \genblk2.pcpi_div_lte_2493_16_n_27 ,
       \genblk2.pcpi_div_lte_2493_16_n_28 ,
       \genblk2.pcpi_div_lte_2493_16_n_29 ;
  wire \genblk2.pcpi_div_lte_2493_16_n_30 ,
       \genblk2.pcpi_div_lte_2493_16_n_31 ,
       \genblk2.pcpi_div_lte_2493_16_n_32 ,
       \genblk2.pcpi_div_lte_2493_16_n_33 ,
       \genblk2.pcpi_div_lte_2493_16_n_34 ,
       \genblk2.pcpi_div_lte_2493_16_n_35 ,
       \genblk2.pcpi_div_lte_2493_16_n_36 ,
       \genblk2.pcpi_div_lte_2493_16_n_37 ;
  wire \genblk2.pcpi_div_lte_2493_16_n_38 ,
       \genblk2.pcpi_div_lte_2493_16_n_39 ,
       \genblk2.pcpi_div_lte_2493_16_n_40 ,
       \genblk2.pcpi_div_lte_2493_16_n_41 ,
       \genblk2.pcpi_div_lte_2493_16_n_42 ,
       \genblk2.pcpi_div_lte_2493_16_n_43 ,
       \genblk2.pcpi_div_lte_2493_16_n_44 ,
       \genblk2.pcpi_div_lte_2493_16_n_45 ;
  wire \genblk2.pcpi_div_lte_2493_16_n_46 ,
       \genblk2.pcpi_div_lte_2493_16_n_47 ,
       \genblk2.pcpi_div_lte_2493_16_n_48 ,
       \genblk2.pcpi_div_lte_2493_16_n_49 ,
       \genblk2.pcpi_div_lte_2493_16_n_50 ,
       \genblk2.pcpi_div_lte_2493_16_n_51 ,
       \genblk2.pcpi_div_lte_2493_16_n_52 ,
       \genblk2.pcpi_div_lte_2493_16_n_53 ;
  wire \genblk2.pcpi_div_lte_2493_16_n_54 ,
       \genblk2.pcpi_div_lte_2493_16_n_55 ,
       \genblk2.pcpi_div_lte_2493_16_n_56 ,
       \genblk2.pcpi_div_lte_2493_16_n_57 ,
       \genblk2.pcpi_div_lte_2493_16_n_58 ,
       \genblk2.pcpi_div_lte_2493_16_n_59 ,
       \genblk2.pcpi_div_lte_2493_16_n_60 ,
       \genblk2.pcpi_div_lte_2493_16_n_61 ;
  wire \genblk2.pcpi_div_lte_2493_16_n_62 ,
       \genblk2.pcpi_div_lte_2493_16_n_63 ,
       \genblk2.pcpi_div_lte_2493_16_n_64 ,
       \genblk2.pcpi_div_lte_2493_16_n_65 ,
       \genblk2.pcpi_div_lte_2493_16_n_66 ,
       \genblk2.pcpi_div_lte_2493_16_n_67 ,
       \genblk2.pcpi_div_lte_2493_16_n_68 ,
       \genblk2.pcpi_div_lte_2493_16_n_69 ;
  wire \genblk2.pcpi_div_lte_2493_16_n_70 ,
       \genblk2.pcpi_div_lte_2493_16_n_71 ,
       \genblk2.pcpi_div_lte_2493_16_n_72 ,
       \genblk2.pcpi_div_lte_2493_16_n_73 ,
       \genblk2.pcpi_div_lte_2493_16_n_74 ,
       \genblk2.pcpi_div_lte_2493_16_n_75 ,
       \genblk2.pcpi_div_lte_2493_16_n_76 ,
       \genblk2.pcpi_div_lte_2493_16_n_77 ;
  wire \genblk2.pcpi_div_lte_2493_16_n_78 ,
       \genblk2.pcpi_div_lte_2493_16_n_79 ,
       \genblk2.pcpi_div_lte_2493_16_n_80 ,
       \genblk2.pcpi_div_lte_2493_16_n_81 ,
       \genblk2.pcpi_div_lte_2493_16_n_82 ,
       \genblk2.pcpi_div_lte_2493_16_n_83 ,
       \genblk2.pcpi_div_lte_2493_16_n_84 ,
       \genblk2.pcpi_div_lte_2493_16_n_85 ;
  wire \genblk2.pcpi_div_lte_2493_16_n_86 ,
       \genblk2.pcpi_div_lte_2493_16_n_87 ,
       \genblk2.pcpi_div_lte_2493_16_n_88 ,
       \genblk2.pcpi_div_lte_2493_16_n_89 ,
       \genblk2.pcpi_div_lte_2493_16_n_90 ,
       \genblk2.pcpi_div_lte_2493_16_n_91 ,
       \genblk2.pcpi_div_lte_2493_16_n_92 ,
       \genblk2.pcpi_div_lte_2493_16_n_93 ;
  wire \genblk2.pcpi_div_lte_2493_16_n_94 ,
       \genblk2.pcpi_div_lte_2493_16_n_95 ,
       \genblk2.pcpi_div_lte_2493_16_n_96 ,
       \genblk2.pcpi_div_lte_2493_16_n_97 ,
       \genblk2.pcpi_div_lte_2493_16_n_98 ,
       \genblk2.pcpi_div_lte_2493_16_n_99 ,
       \genblk2.pcpi_div_lte_2493_16_n_100 ,
       \genblk2.pcpi_div_lte_2493_16_n_101 ;
  wire \genblk2.pcpi_div_lte_2493_16_n_102 ,
       \genblk2.pcpi_div_minus_2470_59_n_324 ,
       \genblk2.pcpi_div_minus_2470_59_n_329 ,
       \genblk2.pcpi_div_minus_2470_59_n_330 ,
       \genblk2.pcpi_div_minus_2470_59_n_335 ,
       \genblk2.pcpi_div_minus_2470_59_n_340 ,
       \genblk2.pcpi_div_minus_2470_59_n_345 ,
       \genblk2.pcpi_div_minus_2470_59_n_350 ;
  wire \genblk2.pcpi_div_minus_2470_59_n_355 ,
       \genblk2.pcpi_div_minus_2470_59_n_360 ,
       \genblk2.pcpi_div_minus_2470_59_n_365 ,
       \genblk2.pcpi_div_minus_2470_59_n_370 ,
       \genblk2.pcpi_div_minus_2470_59_n_375 ,
       \genblk2.pcpi_div_minus_2470_59_n_380 ,
       \genblk2.pcpi_div_minus_2470_59_n_385 ,
       \genblk2.pcpi_div_minus_2470_59_n_390 ;
  wire \genblk2.pcpi_div_minus_2470_59_n_395 ,
       \genblk2.pcpi_div_minus_2470_59_n_400 ,
       \genblk2.pcpi_div_minus_2470_59_n_405 ,
       \genblk2.pcpi_div_minus_2470_59_n_410 ,
       \genblk2.pcpi_div_minus_2470_59_n_415 ,
       \genblk2.pcpi_div_minus_2470_59_n_420 ,
       \genblk2.pcpi_div_minus_2470_59_n_425 ,
       \genblk2.pcpi_div_minus_2470_59_n_430 ;
  wire \genblk2.pcpi_div_minus_2470_59_n_435 ,
       \genblk2.pcpi_div_minus_2470_59_n_440 ,
       \genblk2.pcpi_div_minus_2470_59_n_445 ,
       \genblk2.pcpi_div_minus_2470_59_n_450 ,
       \genblk2.pcpi_div_minus_2470_59_n_455 ,
       \genblk2.pcpi_div_minus_2470_59_n_460 ,
       \genblk2.pcpi_div_minus_2470_59_n_465 ,
       \genblk2.pcpi_div_minus_2470_59_n_470 ;
  wire \genblk2.pcpi_div_minus_2470_59_n_474 ,
       \genblk2.pcpi_div_minus_2470_59_n_476 ,
       \genblk2.pcpi_div_minus_2470_59_n_477 ,
       \genblk2.pcpi_div_minus_2470_59_n_479 ,
       \genblk2.pcpi_div_minus_2470_59_n_481 ,
       \genblk2.pcpi_div_minus_2470_59_n_483 ,
       \genblk2.pcpi_div_minus_2470_59_n_485 ,
       \genblk2.pcpi_div_minus_2470_59_n_487 ;
  wire \genblk2.pcpi_div_minus_2470_59_n_488 ,
       \genblk2.pcpi_div_minus_2470_59_n_492 ,
       \genblk2.pcpi_div_minus_2470_59_n_498 ,
       \genblk2.pcpi_div_minus_2470_59_n_499 ,
       \genblk2.pcpi_div_minus_2470_59_n_500 ,
       \genblk2.pcpi_div_minus_2470_59_n_502 ,
       \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_323 ,
       \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_328 ;
  wire \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_329 ,
       \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_334 ,
       \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_339 ,
       \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_344 ,
       \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_349 ,
       \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_354 ,
       \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_359 ,
       \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_364 ;
  wire \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_369 ,
       \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_374 ,
       \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_379 ,
       \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_384 ,
       \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_389 ,
       \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_394 ,
       \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_399 ,
       \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_404 ;
  wire \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_409 ,
       \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_414 ,
       \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_419 ,
       \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_424 ,
       \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_429 ,
       \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_434 ,
       \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_439 ,
       \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_444 ;
  wire \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_449 ,
       \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_454 ,
       \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_459 ,
       \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_464 ,
       \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_469 ,
       \genblk2.pcpi_div_n_314 , \genblk2.pcpi_div_n_578 ,
       \genblk2.pcpi_div_n_1867 ;
  wire \genblk2.pcpi_div_n_1868 , \genblk2.pcpi_div_n_1869 ,
       \genblk2.pcpi_div_n_1870 , \genblk2.pcpi_div_n_1871 ,
       \genblk2.pcpi_div_n_1872 , \genblk2.pcpi_div_n_1873 ,
       \genblk2.pcpi_div_n_1874 , \genblk2.pcpi_div_n_1875 ;
  wire \genblk2.pcpi_div_n_1876 , \genblk2.pcpi_div_n_1877 ,
       \genblk2.pcpi_div_n_1878 , \genblk2.pcpi_div_n_1879 ,
       \genblk2.pcpi_div_n_1880 , \genblk2.pcpi_div_n_1881 ,
       \genblk2.pcpi_div_n_1882 , \genblk2.pcpi_div_n_1883 ;
  wire \genblk2.pcpi_div_n_1884 , \genblk2.pcpi_div_n_1885 ,
       \genblk2.pcpi_div_n_1886 , \genblk2.pcpi_div_n_1887 ,
       \genblk2.pcpi_div_n_1888 , \genblk2.pcpi_div_n_1889 ,
       \genblk2.pcpi_div_n_1890 , \genblk2.pcpi_div_n_1891 ;
  wire \genblk2.pcpi_div_n_1892 , \genblk2.pcpi_div_n_1893 ,
       \genblk2.pcpi_div_n_1894 , \genblk2.pcpi_div_n_1895 ,
       \genblk2.pcpi_div_n_1896 , \genblk2.pcpi_div_n_1897 ,
       \genblk2.pcpi_div_n_1929 , \genblk2.pcpi_div_n_1930 ;
  wire \genblk2.pcpi_div_n_1931 , \genblk2.pcpi_div_n_1932 ,
       \genblk2.pcpi_div_n_1933 , \genblk2.pcpi_div_n_1934 ,
       \genblk2.pcpi_div_n_1935 , \genblk2.pcpi_div_n_1936 ,
       \genblk2.pcpi_div_n_1937 , \genblk2.pcpi_div_n_1938 ;
  wire \genblk2.pcpi_div_n_1939 , \genblk2.pcpi_div_n_1940 ,
       \genblk2.pcpi_div_n_1941 , \genblk2.pcpi_div_n_1942 ,
       \genblk2.pcpi_div_n_1943 , \genblk2.pcpi_div_n_1944 ,
       \genblk2.pcpi_div_n_1945 , \genblk2.pcpi_div_n_1946 ;
  wire \genblk2.pcpi_div_n_1947 , \genblk2.pcpi_div_n_1948 ,
       \genblk2.pcpi_div_n_1949 , \genblk2.pcpi_div_n_1950 ,
       \genblk2.pcpi_div_n_1951 , \genblk2.pcpi_div_n_1952 ,
       \genblk2.pcpi_div_n_1953 , \genblk2.pcpi_div_n_1954 ;
  wire \genblk2.pcpi_div_n_1955 , \genblk2.pcpi_div_n_1956 ,
       \genblk2.pcpi_div_n_1957 , \genblk2.pcpi_div_n_1958 ,
       \genblk2.pcpi_div_n_1959 , \genblk2.pcpi_div_n_1960 ,
       \genblk2.pcpi_div_n_1961 , \genblk2.pcpi_div_n_1998 ;
  wire \genblk2.pcpi_div_n_1999 , \genblk2.pcpi_div_n_2000 ,
       \genblk2.pcpi_div_n_2001 , \genblk2.pcpi_div_n_2002 ,
       \genblk2.pcpi_div_n_2003 , \genblk2.pcpi_div_n_2004 ,
       \genblk2.pcpi_div_n_2005 , \genblk2.pcpi_div_n_2006 ;
  wire \genblk2.pcpi_div_n_2007 , \genblk2.pcpi_div_n_2008 ,
       \genblk2.pcpi_div_n_2009 , \genblk2.pcpi_div_n_2010 ,
       \genblk2.pcpi_div_n_2011 , \genblk2.pcpi_div_n_2012 ,
       \genblk2.pcpi_div_n_2013 , \genblk2.pcpi_div_n_2014 ;
  wire \genblk2.pcpi_div_n_2015 , \genblk2.pcpi_div_n_2016 ,
       \genblk2.pcpi_div_n_2017 , \genblk2.pcpi_div_n_2018 ,
       \genblk2.pcpi_div_n_2019 , \genblk2.pcpi_div_n_2020 ,
       \genblk2.pcpi_div_n_2021 , \genblk2.pcpi_div_n_2022 ;
  wire \genblk2.pcpi_div_n_2023 , \genblk2.pcpi_div_n_2024 ,
       \genblk2.pcpi_div_n_2025 , \genblk2.pcpi_div_n_2026 ,
       \genblk2.pcpi_div_n_2027 , \genblk2.pcpi_div_n_2028 ,
       \genblk2.pcpi_div_n_2109 , \genblk2.pcpi_div_n_2110 ;
  wire \genblk2.pcpi_div_n_2111 , \genblk2.pcpi_div_n_2112 ,
       \genblk2.pcpi_div_n_2114 , \genblk2.pcpi_div_n_2116 ,
       \genblk2.pcpi_div_n_2118 , \genblk2.pcpi_div_n_2120 ,
       \genblk2.pcpi_div_n_2122 , \genblk2.pcpi_div_n_2124 ;
  wire \genblk2.pcpi_div_n_2126 , \genblk2.pcpi_div_n_2128 ,
       \genblk2.pcpi_div_n_2130 , \genblk2.pcpi_div_n_2132 ,
       \genblk2.pcpi_div_n_2134 , \genblk2.pcpi_div_n_2136 ,
       \genblk2.pcpi_div_n_2138 , \genblk2.pcpi_div_n_2140 ;
  wire \genblk2.pcpi_div_n_2142 , \genblk2.pcpi_div_n_2143 ,
       \genblk2.pcpi_div_n_2144 , \genblk2.pcpi_div_n_2145 ,
       \genblk2.pcpi_div_n_2146 , \genblk2.pcpi_div_n_2147 ,
       \genblk2.pcpi_div_n_2148 , \genblk2.pcpi_div_n_2149 ;
  wire \genblk2.pcpi_div_n_2150 , \genblk2.pcpi_div_n_2151 ,
       \genblk2.pcpi_div_n_2152 , \genblk2.pcpi_div_n_2153 ,
       \genblk2.pcpi_div_n_2154 , \genblk2.pcpi_div_n_2155 ,
       \genblk2.pcpi_div_n_2156 , \genblk2.pcpi_div_n_2157 ;
  wire \genblk2.pcpi_div_n_2158 , \genblk2.pcpi_div_n_2159 ,
       \genblk2.pcpi_div_n_2160 , \genblk2.pcpi_div_n_2161 ,
       \genblk2.pcpi_div_n_2162 , \genblk2.pcpi_div_n_2163 ,
       \genblk2.pcpi_div_n_2164 , \genblk2.pcpi_div_n_2165 ;
  wire \genblk2.pcpi_div_n_2166 , \genblk2.pcpi_div_n_2167 ,
       \genblk2.pcpi_div_n_2168 , \genblk2.pcpi_div_n_2169 ,
       \genblk2.pcpi_div_n_2170 , \genblk2.pcpi_div_n_2171 ,
       \genblk2.pcpi_div_n_2172 , \genblk2.pcpi_div_n_4742 ;
  wire \genblk2.pcpi_div_outsign , \genblk2.pcpi_div_pcpi_wait_q ,
       \genblk2.pcpi_div_running ,
       \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1132 ,
       \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1134 ,
       \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1136 ,
       \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1138 ,
       \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1140 ;
  wire \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1142 ,
       \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1144 ,
       \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1146 ,
       \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1148 ,
       \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1150 ,
       \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1152 ,
       \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1154 ,
       \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1156 ;
  wire \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1158 ,
       \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1160 ,
       \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1162 ,
       \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1164 ,
       \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1166 ,
       \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1168 ,
       \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1170 ,
       \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1172 ;
  wire \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1174 ,
       \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1176 ,
       \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1178 ,
       \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1180 ,
       \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1182 ,
       \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1184 ,
       \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1186 ,
       \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1188 ;
  wire \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1190 ,
       \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1194 ,
       \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1213 ,
       inc_add_382_74_n_207, inc_add_382_74_n_212,
       inc_add_382_74_n_217, inc_add_382_74_n_222, inc_add_382_74_n_227;
  wire inc_add_382_74_n_232, inc_add_382_74_n_237,
       inc_add_382_74_n_242, inc_add_382_74_n_247,
       inc_add_382_74_n_252, inc_add_382_74_n_257,
       inc_add_382_74_n_262, inc_add_382_74_n_267;
  wire inc_add_382_74_n_272, inc_add_382_74_n_277,
       inc_add_382_74_n_282, inc_add_382_74_n_287,
       inc_add_382_74_n_292, inc_add_382_74_n_297,
       inc_add_382_74_n_302, inc_add_382_74_n_305;
  wire inc_add_382_74_n_309, inc_add_382_74_n_314,
       inc_add_382_74_n_319, inc_add_382_74_n_324,
       inc_add_382_74_n_329, inc_add_382_74_n_332,
       inc_add_382_74_n_336, inc_add_382_74_n_341;
  wire inc_add_1428_40_n_445, inc_add_1428_40_n_450,
       inc_add_1428_40_n_455, inc_add_1428_40_n_460,
       inc_add_1428_40_n_465, inc_add_1428_40_n_470,
       inc_add_1428_40_n_475, inc_add_1428_40_n_480;
  wire inc_add_1428_40_n_485, inc_add_1428_40_n_490,
       inc_add_1428_40_n_495, inc_add_1428_40_n_500,
       inc_add_1428_40_n_505, inc_add_1428_40_n_510,
       inc_add_1428_40_n_515, inc_add_1428_40_n_520;
  wire inc_add_1428_40_n_525, inc_add_1428_40_n_530,
       inc_add_1428_40_n_535, inc_add_1428_40_n_540,
       inc_add_1428_40_n_545, inc_add_1428_40_n_550,
       inc_add_1428_40_n_555, inc_add_1428_40_n_560;
  wire inc_add_1428_40_n_565, inc_add_1428_40_n_570,
       inc_add_1428_40_n_575, inc_add_1428_40_n_580,
       inc_add_1428_40_n_585, inc_add_1428_40_n_590,
       inc_add_1428_40_n_595, inc_add_1428_40_n_600;
  wire inc_add_1428_40_n_605, inc_add_1428_40_n_610,
       inc_add_1428_40_n_615, inc_add_1428_40_n_620,
       inc_add_1428_40_n_625, inc_add_1428_40_n_630,
       inc_add_1428_40_n_635, inc_add_1428_40_n_640;
  wire inc_add_1428_40_n_645, inc_add_1428_40_n_650,
       inc_add_1428_40_n_655, inc_add_1428_40_n_660,
       inc_add_1428_40_n_665, inc_add_1428_40_n_670,
       inc_add_1428_40_n_675, inc_add_1428_40_n_680;
  wire inc_add_1428_40_n_685, inc_add_1428_40_n_688,
       inc_add_1428_40_n_692, inc_add_1428_40_n_695,
       inc_add_1428_40_n_699, inc_add_1428_40_n_704,
       inc_add_1428_40_n_709, inc_add_1428_40_n_714;
  wire inc_add_1428_40_n_719, inc_add_1428_40_n_722,
       inc_add_1428_40_n_726, inc_add_1428_40_n_731,
       inc_add_1428_40_n_736, inc_add_1428_40_n_741,
       inc_add_1559_34_n_445, inc_add_1559_34_n_450;
  wire inc_add_1559_34_n_455, inc_add_1559_34_n_460,
       inc_add_1559_34_n_465, inc_add_1559_34_n_470,
       inc_add_1559_34_n_475, inc_add_1559_34_n_480,
       inc_add_1559_34_n_485, inc_add_1559_34_n_490;
  wire inc_add_1559_34_n_495, inc_add_1559_34_n_500,
       inc_add_1559_34_n_505, inc_add_1559_34_n_510,
       inc_add_1559_34_n_515, inc_add_1559_34_n_520,
       inc_add_1559_34_n_525, inc_add_1559_34_n_530;
  wire inc_add_1559_34_n_535, inc_add_1559_34_n_540,
       inc_add_1559_34_n_545, inc_add_1559_34_n_550,
       inc_add_1559_34_n_555, inc_add_1559_34_n_560,
       inc_add_1559_34_n_565, inc_add_1559_34_n_570;
  wire inc_add_1559_34_n_575, inc_add_1559_34_n_580,
       inc_add_1559_34_n_585, inc_add_1559_34_n_590,
       inc_add_1559_34_n_595, inc_add_1559_34_n_600,
       inc_add_1559_34_n_605, inc_add_1559_34_n_610;
  wire inc_add_1559_34_n_615, inc_add_1559_34_n_620,
       inc_add_1559_34_n_625, inc_add_1559_34_n_630,
       inc_add_1559_34_n_635, inc_add_1559_34_n_640,
       inc_add_1559_34_n_645, inc_add_1559_34_n_650;
  wire inc_add_1559_34_n_655, inc_add_1559_34_n_660,
       inc_add_1559_34_n_665, inc_add_1559_34_n_670,
       inc_add_1559_34_n_675, inc_add_1559_34_n_680,
       inc_add_1559_34_n_685, inc_add_1559_34_n_688;
  wire inc_add_1559_34_n_692, inc_add_1559_34_n_695,
       inc_add_1559_34_n_699, inc_add_1559_34_n_704,
       inc_add_1559_34_n_709, inc_add_1559_34_n_714,
       inc_add_1559_34_n_719, inc_add_1559_34_n_722;
  wire inc_add_1559_34_n_726, inc_add_1559_34_n_731,
       inc_add_1559_34_n_736, inc_add_1559_34_n_741, instr_add,
       instr_addi, instr_and, instr_andi;
  wire instr_auipc, instr_beq, instr_bge, instr_bgeu, instr_blt,
       instr_bltu, instr_bne, instr_ecall_ebreak;
  wire instr_jal, instr_jalr, instr_lb, instr_lbu, instr_lh, instr_lhu,
       instr_lui, instr_lw;
  wire instr_or, instr_ori, instr_rdcycle, instr_rdcycleh,
       instr_rdinstr, instr_rdinstrh, instr_sb, instr_sh;
  wire instr_sll, instr_slli, instr_slt, instr_slti, instr_sltiu,
       instr_sltu, instr_sra, instr_srai;
  wire instr_srl, instr_srli, instr_sub, instr_sw, instr_xor,
       instr_xori, is_alu_reg_imm, is_alu_reg_reg;
  wire is_beq_bne_blt_bge_bltu_bgeu, is_compare,
       is_jalr_addi_slti_sltiu_xori_ori_andi, is_lb_lh_lw_lbu_lhu,
       is_lbu_lhu_lw, is_lui_auipc_jal,
       is_lui_auipc_jal_jalr_addi_add_sub, is_sb_sh_sw;
  wire is_sll_srl_sra, is_slli_srli_srai, is_slti_blt_slt,
       is_sltiu_bltu_sltu, last_mem_valid, latched_branch,
       latched_compr, latched_is_lb;
  wire latched_is_lh, latched_is_lu, latched_stalu, latched_store,
       mem_do_prefetch, mem_do_rdata, mem_do_rinst, mem_do_wdata;
  wire mem_done, mem_la_firstword_reg, mem_la_firstword_xfer,
       mem_la_secondword, mem_valid_9465, mem_xfer, n_0, n_1;
  wire n_2, n_3, n_4, n_5, n_6, n_7, n_8, n_9;
  wire n_10, n_11, n_12, n_13, n_14, n_15, n_16, n_17;
  wire n_18, n_19, n_20, n_21, n_22, n_23, n_24, n_25;
  wire n_26, n_27, n_28, n_29, n_30, n_31, n_32, n_33;
  wire n_34, n_35, n_36, n_37, n_38, n_39, n_40, n_42;
  wire n_46, n_48, n_50, n_52, n_54, n_56, n_60, n_62;
  wire n_64, n_66, n_68, n_70, n_72, n_74, n_76, n_78;
  wire n_80, n_82, n_84, n_86, n_88, n_90, n_92, n_94;
  wire n_96, n_98, n_100, n_102, n_104, n_106, n_108, n_110;
  wire n_112, n_113, n_114, n_115, n_119, n_120, n_122, n_130;
  wire n_136, n_138, n_142, n_144, n_146, n_150, n_152, n_154;
  wire n_156, n_158, n_160, n_162, n_164, n_166, n_168, n_170;
  wire n_172, n_174, n_176, n_178, n_180, n_182, n_184, n_186;
  wire n_188, n_190, n_192, n_194, n_196, n_198, n_200, n_202;
  wire n_204, n_206, n_208, n_210, n_212, n_214, n_216, n_218;
  wire n_219, n_222, n_228, n_258, n_268, n_276, n_277, n_278;
  wire n_279, n_283, n_288, n_289, n_290, n_291, n_293, n_294;
  wire n_296, n_297, n_300, n_301, n_302, n_303, n_305, n_306;
  wire n_307, n_308, n_309, n_310, n_311, n_313, n_314, n_316;
  wire n_317, n_318, n_320, n_321, n_323, n_324, n_325, n_326;
  wire n_327, n_329, n_331, n_332, n_333, n_334, n_335, n_338;
  wire n_340, n_341, n_342, n_343, n_344, n_345, n_347, n_348;
  wire n_349, n_353, n_355, n_356, n_358, n_360, n_362, n_364;
  wire n_366, n_368, n_370, n_372, n_374, n_376, n_378, n_380;
  wire n_382, n_384, n_386, n_388, n_390, n_392, n_394, n_396;
  wire n_398, n_400, n_402, n_404, n_406, n_408, n_412, n_414;
  wire n_416, n_418, n_419, n_421, n_423, n_424, n_425, n_427;
  wire n_429, n_431, n_432, n_434, n_436, n_437, n_438, n_439;
  wire n_440, n_441, n_442, n_444, n_445, n_446, n_448, n_450;
  wire n_452, n_454, n_456, n_458, n_460, n_462, n_464, n_466;
  wire n_468, n_470, n_472, n_474, n_476, n_478, n_480, n_482;
  wire n_484, n_486, n_488, n_490, n_492, n_494, n_496, n_498;
  wire n_500, n_502, n_503, n_504, n_505, n_506, n_508, n_510;
  wire n_512, n_514, n_516, n_518, n_520, n_522, n_524, n_526;
  wire n_528, n_530, n_532, n_534, n_536, n_537, n_538, n_540;
  wire n_542, n_543, n_544, n_545, n_547, n_548, n_550, n_552;
  wire n_555, n_558, n_562, n_564, n_565, n_567, n_572, n_573;
  wire n_574, n_576, n_577, n_578, n_579, n_580, n_581, n_582;
  wire n_583, n_586, n_587, n_588, n_589, n_590, n_591, n_592;
  wire n_593, n_594, n_595, n_596, n_597, n_598, n_599, n_600;
  wire n_601, n_602, n_603, n_604, n_605, n_606, n_607, n_608;
  wire n_609, n_611, n_613, n_615, n_616, n_619, n_622, n_624;
  wire n_625, n_627, n_628, n_629, n_630, n_633, n_634, n_635;
  wire n_636, n_637, n_638, n_639, n_640, n_641, n_642, n_643;
  wire n_644, n_645, n_646, n_647, n_648, n_649, n_650, n_651;
  wire n_652, n_653, n_654, n_655, n_656, n_657, n_658, n_659;
  wire n_662, n_663, n_664, n_665, n_666, n_667, n_668, n_671;
  wire n_672, n_673, n_674, n_675, n_676, n_677, n_678, n_679;
  wire n_680, n_681, n_682, n_683, n_685, n_686, n_687, n_688;
  wire n_689, n_690, n_691, n_692, n_693, n_695, n_696, n_697;
  wire n_702, n_703, n_704, n_705, n_706, n_707, n_709, n_712;
  wire n_713, n_714, n_715, n_716, n_717, n_718, n_721, n_722;
  wire n_723, n_725, n_726, n_727, n_728, n_729, n_730, n_731;
  wire n_732, n_733, n_734, n_735, n_736, n_739, n_740, n_744;
  wire n_745, n_746, n_747, n_751, n_752, n_756, n_759, n_760;
  wire n_761, n_762, n_763, n_764, n_765, n_766, n_767, n_768;
  wire n_769, n_770, n_771, n_772, n_773, n_774, n_775, n_776;
  wire n_777, n_778, n_779, n_781, n_782, n_783, n_784, n_785;
  wire n_786, n_787, n_788, n_789, n_790, n_791, n_792, n_793;
  wire n_794, n_795, n_796, n_797, n_798, n_799, n_800, n_801;
  wire n_802, n_803, n_804, n_805, n_806, n_807, n_808, n_809;
  wire n_810, n_811, n_812, n_813, n_814, n_815, n_816, n_817;
  wire n_818, n_819, n_820, n_821, n_822, n_823, n_824, n_825;
  wire n_826, n_827, n_828, n_829, n_830, n_832, n_833, n_839;
  wire n_842, n_843, n_844, n_845, n_846, n_847, n_848, n_849;
  wire n_850, n_851, n_852, n_853, n_854, n_855, n_856, n_857;
  wire n_858, n_859, n_860, n_861, n_862, n_863, n_865, n_866;
  wire n_867, n_868, n_869, n_870, n_871, n_873, n_874, n_875;
  wire n_876, n_877, n_878, n_879, n_880, n_881, n_882, n_883;
  wire n_884, n_885, n_886, n_887, n_888, n_889, n_890, n_891;
  wire n_892, n_893, n_894, n_895, n_896, n_897, n_898, n_899;
  wire n_900, n_901, n_902, n_903, n_904, n_905, n_906, n_907;
  wire n_908, n_909, n_910, n_911, n_912, n_913, n_914, n_915;
  wire n_916, n_917, n_918, n_919, n_920, n_921, n_922, n_923;
  wire n_924, n_925, n_926, n_927, n_928, n_929, n_930, n_931;
  wire n_932, n_933, n_934, n_935, n_936, n_937, n_938, n_939;
  wire n_940, n_941, n_942, n_943, n_944, n_945, n_946, n_947;
  wire n_948, n_949, n_950, n_951, n_952, n_953, n_954, n_957;
  wire n_960, n_961, n_962, n_963, n_964, n_965, n_966, n_967;
  wire n_968, n_969, n_970, n_971, n_972, n_973, n_974, n_975;
  wire n_976, n_977, n_978, n_979, n_980, n_981, n_982, n_983;
  wire n_984, n_985, n_986, n_987, n_988, n_989, n_990, n_991;
  wire n_992, n_993, n_994, n_995, n_996, n_997, n_998, n_999;
  wire n_1000, n_1001, n_1002, n_1003, n_1004, n_1005, n_1006, n_1007;
  wire n_1008, n_1009, n_1010, n_1011, n_1012, n_1013, n_1014, n_1015;
  wire n_1016, n_1017, n_1018, n_1019, n_1020, n_1021, n_1022, n_1023;
  wire n_1024, n_1025, n_1026, n_1027, n_1028, n_1029, n_1030, n_1031;
  wire n_1032, n_1033, n_1034, n_1035, n_1036, n_1037, n_1038, n_1039;
  wire n_1040, n_1041, n_1042, n_1043, n_1044, n_1045, n_1046, n_1047;
  wire n_1048, n_1049, n_1050, n_1051, n_1052, n_1053, n_1054, n_1055;
  wire n_1056, n_1057, n_1058, n_1059, n_1060, n_1061, n_1062, n_1063;
  wire n_1064, n_1065, n_1066, n_1067, n_1068, n_1069, n_1070, n_1071;
  wire n_1072, n_1073, n_1074, n_1075, n_1076, n_1077, n_1078, n_1079;
  wire n_1080, n_1081, n_1082, n_1083, n_1084, n_1085, n_1086, n_1087;
  wire n_1088, n_1089, n_1090, n_1091, n_1092, n_1093, n_1094, n_1095;
  wire n_1096, n_1097, n_1098, n_1099, n_1100, n_1101, n_1102, n_1103;
  wire n_1104, n_1105, n_1106, n_1107, n_1108, n_1109, n_1110, n_1111;
  wire n_1112, n_1113, n_1114, n_1115, n_1116, n_1117, n_1118, n_1119;
  wire n_1120, n_1121, n_1122, n_1123, n_1124, n_1125, n_1126, n_1127;
  wire n_1128, n_1129, n_1130, n_1131, n_1132, n_1133, n_1134, n_1135;
  wire n_1136, n_1137, n_1138, n_1139, n_1140, n_1141, n_1142, n_1143;
  wire n_1144, n_1145, n_1146, n_1147, n_1148, n_1149, n_1150, n_1151;
  wire n_1152, n_1153, n_1154, n_1155, n_1156, n_1157, n_1158, n_1159;
  wire n_1160, n_1161, n_1162, n_1165, n_1166, n_1167, n_1168, n_1169;
  wire n_1170, n_1173, n_1174, n_1176, n_1177, n_1178, n_1181, n_1182;
  wire n_1183, n_1184, n_1185, n_1186, n_1187, n_1188, n_1190, n_1191;
  wire n_1192, n_1193, n_1194, n_1195, n_1196, n_1197, n_1198, n_1199;
  wire n_1200, n_1201, n_1202, n_1203, n_1204, n_1205, n_1206, n_1207;
  wire n_1208, n_1209, n_1210, n_1211, n_1212, n_1213, n_1214, n_1215;
  wire n_1216, n_1231, n_1232, n_1233, n_1234, n_1248, n_1254, n_1256;
  wire n_1258, n_1259, n_1261, n_1263, n_1266, n_1267, n_1269, n_1271;
  wire n_1272, n_1278, n_1280, n_1281, n_1282, n_1299, n_1300, n_1301;
  wire n_1302, n_1303, n_1304, n_1305, n_1306, n_1307, n_1308, n_1310;
  wire n_1318, n_1319, n_1320, n_1321, n_1322, n_1323, n_1324, n_1325;
  wire n_1326, n_1327, n_1328, n_1329, n_1330, n_1331, n_1332, n_1333;
  wire n_1334, n_1335, n_1336, n_1337, n_1338, n_1339, n_1340, n_1341;
  wire n_1342, n_1343, n_1344, n_1345, n_1346, n_1347, n_1348, n_1349;
  wire n_1350, n_1351, n_1352, n_1353, n_1354, n_1355, n_1356, n_1357;
  wire n_1358, n_1359, n_1360, n_1361, n_1362, n_1363, n_1364, n_1365;
  wire n_1366, n_1367, n_1368, n_1369, n_1370, n_1372, n_1373, n_1374;
  wire n_1375, n_1376, n_1377, n_1378, n_1379, n_1380, n_1381, n_1382;
  wire n_1383, n_1384, n_1385, n_1386, n_1387, n_1388, n_1389, n_1390;
  wire n_1391, n_1392, n_1393, n_1394, n_1395, n_1396, n_1397, n_1398;
  wire n_1399, n_1400, n_1401, n_1402, n_1403, n_1404, n_1405, n_1406;
  wire n_1407, n_1408, n_1409, n_1410, n_1411, n_1412, n_1413, n_1414;
  wire n_1415, n_1416, n_1417, n_1418, n_1419, n_1420, n_1421, n_1422;
  wire n_1423, n_1424, n_1425, n_1426, n_1427, n_1428, n_1430, n_1431;
  wire n_1432, n_1433, n_1434, n_1435, n_1436, n_1437, n_1438, n_1440;
  wire n_1441, n_1442, n_1443, n_1444, n_1445, n_1446, n_1447, n_1448;
  wire n_1449, n_1451, n_1452, n_1453, n_1454, n_1455, n_1456, n_1457;
  wire n_1458, n_1459, n_1460, n_1461, n_1462, n_1464, n_1465, n_1466;
  wire n_1467, n_1468, n_1469, n_1470, n_1472, n_1473, n_1474, n_1475;
  wire n_1476, n_1477, n_1478, n_1479, n_1480, n_1482, n_1488, n_1512;
  wire n_1513, n_1514, n_1515, n_1517, n_1518, n_1523, n_1525, n_1526;
  wire n_1527, n_1528, n_1529, n_1530, n_1531, n_1532, n_1533, n_1534;
  wire n_1535, n_1536, n_1537, n_1538, n_1539, n_1540, n_1541, n_1542;
  wire n_1543, n_1544, n_1545, n_1546, n_1547, n_1548, n_1549, n_1550;
  wire n_1552, n_1553, n_1554, n_1555, n_1556, n_1557, n_1558, n_1559;
  wire n_1560, n_1584, n_1585, n_1586, n_1588, n_1589, n_1590, n_1591;
  wire n_1592, n_1593, n_1594, n_1595, n_1596, n_1597, n_1598, n_1599;
  wire n_1600, n_1601, n_1602, n_1603, n_1604, n_1605, n_1606, n_1607;
  wire n_1608, n_1609, n_1610, n_1611, n_1613, n_1614, n_1615, n_1616;
  wire n_1617, n_1618, n_1619, n_1620, n_1621, n_1622, n_1623, n_1624;
  wire n_1625, n_1626, n_1627, n_1628, n_1629, n_1630, n_1631, n_1632;
  wire n_1633, n_1634, n_1635, n_1636, n_1637, n_1638, n_1639, n_1640;
  wire n_1654, n_1655, n_1656, n_1657, n_1658, n_1659, n_1660, n_1661;
  wire n_1662, n_1663, n_1664, n_1665, n_1666, n_1667, n_1668, n_1669;
  wire n_1670, n_1671, n_1672, n_1673, n_1674, n_1675, n_1676, n_1677;
  wire n_1678, n_1679, n_1680, n_1681, n_1682, n_1683, n_1684, n_1685;
  wire n_1686, n_1687, n_1688, n_1689, n_1690, n_1691, n_1692, n_1693;
  wire n_1694, n_1695, n_1696, n_1697, n_1698, n_1699, n_1700, n_1701;
  wire n_1702, n_1703, n_1704, n_1705, n_1706, n_1707, n_1708, n_1710;
  wire n_1711, n_1712, n_1713, n_1714, n_1715, n_1716, n_1717, n_1718;
  wire n_1719, n_1720, n_1721, n_1722, n_1723, n_1724, n_1725, n_1726;
  wire n_1727, n_1728, n_1729, n_1730, n_1731, n_1732, n_1733, n_1734;
  wire n_1735, n_1736, n_1737, n_1738, n_1739, n_1742, n_1743, n_1744;
  wire n_1745, n_1746, n_1755, n_1756, n_1757, n_1758, n_1759, n_1760;
  wire n_1761, n_1762, n_1763, n_1764, n_1765, n_1766, n_1767, n_1768;
  wire n_1769, n_1770, n_1771, n_1772, n_1773, n_1774, n_1775, n_1776;
  wire n_1777, n_1778, n_1779, n_1780, n_1781, n_1782, n_1783, n_1784;
  wire n_1785, n_1786, n_1787, n_1788, n_1789, n_1790, n_1791, n_1792;
  wire n_1793, n_1794, n_1795, n_1796, n_1797, n_1798, n_1799, n_1800;
  wire n_1801, n_1802, n_1803, n_1804, n_1805, n_1806, n_1807, n_1808;
  wire n_1809, n_1810, n_1811, n_1812, n_1813, n_1814, n_1815, n_1816;
  wire n_1817, n_1818, n_1819, n_1820, n_1821, n_1822, n_1823, n_1824;
  wire n_1825, n_1826, n_1827, n_1828, n_1829, n_1830, n_1831, n_1832;
  wire n_1833, n_1834, n_1835, n_1836, n_1837, n_1838, n_1839, n_1840;
  wire n_1841, n_1842, n_1843, n_1844, n_1845, n_1846, n_1847, n_1848;
  wire n_1849, n_1850, n_1851, n_1852, n_1853, n_1854, n_1855, n_1856;
  wire n_1857, n_1858, n_1859, n_1860, n_1861, n_1862, n_1863, n_1864;
  wire n_1865, n_1866, n_1868, n_1869, n_1870, n_1871, n_1872, n_1873;
  wire n_1874, n_1875, n_1876, n_1877, n_1878, n_1879, n_1880, n_1881;
  wire n_1882, n_1883, n_1884, n_1885, n_1886, n_1887, n_1888, n_1889;
  wire n_1890, n_1891, n_1892, n_1893, n_1894, n_1895, n_1896, n_1897;
  wire n_1898, n_1899, n_1900, n_1901, n_1902, n_1903, n_1904, n_1905;
  wire n_1906, n_1907, n_1908, n_1909, n_1910, n_1911, n_1912, n_1913;
  wire n_1914, n_1915, n_1916, n_1917, n_1918, n_1919, n_1920, n_1921;
  wire n_1922, n_1923, n_1924, n_1925, n_1926, n_1927, n_1928, n_1929;
  wire n_1930, n_1931, n_1932, n_1933, n_1934, n_1935, n_1937, n_1938;
  wire n_1939, n_1940, n_1941, n_1943, n_1944, n_1946, n_1947, n_1948;
  wire n_1949, n_1950, n_1951, n_1953, n_1954, n_1955, n_1956, n_1957;
  wire n_1958, n_1974, n_1976, n_1977, n_1979, n_1980, n_1981, n_1982;
  wire n_1983, n_1984, n_1985, n_1986, n_1987, n_1988, n_1989, n_1990;
  wire n_1991, n_1992, n_1993, n_1994, n_1995, n_1996, n_1997, n_2009;
  wire n_2010, n_2011, n_2012, n_2013, n_2014, n_2015, n_2016, n_2017;
  wire n_2018, n_2019, n_2020, n_2021, n_2022, n_2023, n_2024, n_2025;
  wire n_2026, n_2027, n_2028, n_2029, n_2030, n_2031, n_2032, n_2033;
  wire n_2034, n_2035, n_2036, n_2037, n_2038, n_2039, n_2040, n_2041;
  wire n_2042, n_2043, n_2044, n_2045, n_2046, n_2047, n_2048, n_2050;
  wire n_2051, n_2052, n_2053, n_2054, n_2055, n_2056, n_2057, n_2058;
  wire n_2059, n_2060, n_2061, n_2062, n_2063, n_2064, n_2065, n_2066;
  wire n_2067, n_2068, n_2069, n_2070, n_2071, n_2072, n_2073, n_2074;
  wire n_2075, n_2076, n_2077, n_2078, n_2079, n_2080, n_2081, n_2082;
  wire n_2083, n_2084, n_2085, n_2086, n_2087, n_2088, n_2089, n_2090;
  wire n_2091, n_2092, n_2093, n_2094, n_2095, n_2096, n_2097, n_2098;
  wire n_2099, n_2100, n_2101, n_2102, n_2103, n_2104, n_2105, n_2106;
  wire n_2107, n_2108, n_2109, n_2110, n_2111, n_2113, n_2114, n_2115;
  wire n_2116, n_2117, n_2118, n_2119, n_2120, n_2121, n_2122, n_2123;
  wire n_2124, n_2125, n_2126, n_2127, n_2128, n_2131, n_2137, n_2140;
  wire n_2143, n_2144, n_2145, n_2146, n_2150, n_2151, n_2152, n_2153;
  wire n_2154, n_2155, n_2156, n_2157, n_2158, n_2159, n_2161, n_2162;
  wire n_2163, n_2164, n_2165, n_2166, n_2167, n_2168, n_2169, n_2170;
  wire n_2171, n_2172, n_2173, n_2174, n_2175, n_2176, n_2177, n_2178;
  wire n_2179, n_2180, n_2181, n_2182, n_2183, n_2184, n_2185, n_2186;
  wire n_2187, n_2188, n_2189, n_2190, n_2191, n_2192, n_2193, n_2194;
  wire n_2195, n_2196, n_2197, n_2198, n_2199, n_2200, n_2201, n_2202;
  wire n_2203, n_2204, n_2205, n_2206, n_2207, n_2208, n_2209, n_2210;
  wire n_2211, n_2212, n_2213, n_2214, n_2215, n_2216, n_2217, n_2218;
  wire n_2219, n_2220, n_2221, n_2222, n_2223, n_2224, n_2225, n_2226;
  wire n_2227, n_2228, n_2229, n_2230, n_2231, n_2232, n_2233, n_2234;
  wire n_2235, n_2236, n_2237, n_2238, n_2239, n_2240, n_2241, n_2242;
  wire n_2243, n_2244, n_2245, n_2246, n_2247, n_2248, n_2249, n_2250;
  wire n_2251, n_2252, n_2253, n_2254, n_2255, n_2256, n_2257, n_2258;
  wire n_2259, n_2260, n_2261, n_2262, n_2263, n_2264, n_2265, n_2266;
  wire n_2267, n_2268, n_2269, n_2270, n_2271, n_2272, n_2273, n_2274;
  wire n_2275, n_2276, n_2277, n_2278, n_2279, n_2280, n_2281, n_2282;
  wire n_2283, n_2284, n_2285, n_2286, n_2287, n_2288, n_2289, n_2290;
  wire n_2291, n_2292, n_2293, n_2294, n_2295, n_2296, n_2297, n_2298;
  wire n_2299, n_2300, n_2301, n_2302, n_2303, n_2304, n_2305, n_2306;
  wire n_2307, n_2308, n_2309, n_2310, n_2311, n_2312, n_2314, n_2315;
  wire n_2316, n_2317, n_2318, n_2319, n_2320, n_2321, n_2322, n_2323;
  wire n_2324, n_2325, n_2326, n_2327, n_2328, n_2329, n_2330, n_2332;
  wire n_2333, n_2334, n_2335, n_2336, n_2337, n_2338, n_2339, n_2340;
  wire n_2341, n_2342, n_2343, n_2344, n_2345, n_2346, n_2347, n_2348;
  wire n_2349, n_2350, n_2351, n_2352, n_2353, n_2354, n_2355, n_2356;
  wire n_2357, n_2358, n_2359, n_2360, n_2361, n_2362, n_2363, n_2364;
  wire n_2365, n_2366, n_2367, n_2368, n_2369, n_2370, n_2371, n_2372;
  wire n_2377, n_2378, n_2379, n_2380, n_2381, n_2382, n_2383, n_2384;
  wire n_2385, n_2386, n_2387, n_2388, n_2389, n_2390, n_2391, n_2392;
  wire n_2393, n_2394, n_2395, n_2396, n_2397, n_2398, n_2399, n_2400;
  wire n_2401, n_2402, n_2403, n_2404, n_2405, n_2406, n_2407, n_2408;
  wire n_2409, n_2410, n_2411, n_2412, n_2414, n_2415, n_2416, n_2417;
  wire n_2418, n_2421, n_2422, n_2423, n_2424, n_2425, n_2426, n_2427;
  wire n_2428, n_2429, n_2430, n_2431, n_2433, n_2434, n_2435, n_2436;
  wire n_2437, n_2438, n_2439, n_2440, n_2441, n_2442, n_2443, n_2444;
  wire n_2445, n_2446, n_2447, n_2448, n_2449, n_2450, n_2451, n_2452;
  wire n_2453, n_2454, n_2455, n_2456, n_2457, n_2458, n_2459, n_2460;
  wire n_2461, n_2462, n_2463, n_2464, n_2465, n_2466, n_2467, n_2468;
  wire n_2469, n_2470, n_2471, n_2472, n_2473, n_2474, n_2475, n_2476;
  wire n_2477, n_2478, n_2479, n_2480, n_2481, n_2482, n_2483, n_2484;
  wire n_2485, n_2486, n_2487, n_2488, n_2489, n_2490, n_2491, n_2492;
  wire n_2493, n_2494, n_2495, n_2496, n_2497, n_2498, n_2499, n_2500;
  wire n_2502, n_2503, n_2504, n_2505, n_2506, n_2508, n_2509, n_2510;
  wire n_2511, n_2512, n_2513, n_2514, n_2515, n_2516, n_2517, n_2518;
  wire n_2519, n_2520, n_2521, n_2522, n_2523, n_2524, n_2525, n_2526;
  wire n_2527, n_2528, n_2529, n_2530, n_2531, n_2532, n_2533, n_2534;
  wire n_2535, n_2536, n_2537, n_2538, n_2539, n_2540, n_2541, n_2542;
  wire n_2543, n_2544, n_2545, n_2546, n_2547, n_2548, n_2549, n_2550;
  wire n_2551, n_2552, n_2553, n_2554, n_2555, n_2556, n_2557, n_2558;
  wire n_2559, n_2560, n_2561, n_2562, n_2563, n_2564, n_2565, n_2566;
  wire n_2567, n_2568, n_2569, n_2570, n_2571, n_2572, n_2573, n_2574;
  wire n_2575, n_2576, n_2577, n_2578, n_2579, n_2580, n_2581, n_2582;
  wire n_2584, n_2585, n_2586, n_2587, n_2588, n_2589, n_2590, n_2591;
  wire n_2592, n_2593, n_2594, n_2595, n_2597, n_2598, n_2599, n_2600;
  wire n_2601, n_2602, n_2603, n_2604, n_2605, n_2606, n_2607, n_2608;
  wire n_2609, n_2610, n_2611, n_2612, n_2613, n_2614, n_2615, n_2616;
  wire n_2617, n_2618, n_2619, n_2620, n_2621, n_2622, n_2623, n_2624;
  wire n_2625, n_2626, n_2627, n_2628, n_2629, n_2630, n_2631, n_2632;
  wire n_2633, n_2634, n_2635, n_2636, n_2637, n_2638, n_2639, n_2640;
  wire n_2641, n_2642, n_2643, n_2644, n_2645, n_2646, n_2647, n_2648;
  wire n_2649, n_2650, n_2651, n_2652, n_2653, n_2654, n_2655, n_2656;
  wire n_2657, n_2658, n_2659, n_2660, n_2661, n_2662, n_2663, n_2664;
  wire n_2665, n_2666, n_2667, n_2668, n_2669, n_2670, n_2671, n_2672;
  wire n_2673, n_2674, n_2675, n_2676, n_2677, n_2678, n_2679, n_2680;
  wire n_2681, n_2682, n_2683, n_2684, n_2685, n_2686, n_2687, n_2688;
  wire n_2689, n_2690, n_2691, n_2692, n_2693, n_2694, n_2695, n_2696;
  wire n_2697, n_2698, n_2699, n_2700, n_2701, n_2702, n_2703, n_2704;
  wire n_2705, n_2706, n_2707, n_2708, n_2709, n_2710, n_2711, n_2712;
  wire n_2713, n_2714, n_2715, n_2716, n_2717, n_2718, n_2719, n_2720;
  wire n_2721, n_2722, n_2723, n_2724, n_2725, n_2726, n_2727, n_2728;
  wire n_2729, n_2730, n_2731, n_2732, n_2733, n_2734, n_2735, n_2736;
  wire n_2737, n_2738, n_2739, n_2740, n_2741, n_2742, n_2743, n_2744;
  wire n_2745, n_2746, n_2747, n_2748, n_2749, n_2750, n_2751, n_2752;
  wire n_2753, n_2754, n_2755, n_2756, n_2757, n_2758, n_2759, n_2760;
  wire n_2761, n_2762, n_2763, n_2764, n_2765, n_2766, n_2767, n_2768;
  wire n_2769, n_2770, n_2771, n_2772, n_2773, n_2774, n_2775, n_2776;
  wire n_2777, n_2778, n_2779, n_2780, n_2781, n_2782, n_2783, n_2784;
  wire n_2785, n_2786, n_2787, n_2788, n_2789, n_2790, n_2791, n_2792;
  wire n_2793, n_2794, n_2795, n_2796, n_2797, n_2798, n_2799, n_2800;
  wire n_2801, n_2802, n_2803, n_2804, n_2805, n_2806, n_2807, n_2808;
  wire n_2809, n_2810, n_2811, n_2812, n_2813, n_2814, n_2815, n_2816;
  wire n_2817, n_2818, n_2819, n_2820, n_2821, n_2822, n_2823, n_2824;
  wire n_2825, n_2826, n_2827, n_2828, n_2829, n_2830, n_2831, n_2832;
  wire n_2833, n_2834, n_2835, n_2836, n_2837, n_2838, n_2839, n_2840;
  wire n_2841, n_2842, n_2843, n_2844, n_2845, n_2846, n_2847, n_2848;
  wire n_2849, n_2850, n_2851, n_2852, n_2853, n_2854, n_2855, n_2856;
  wire n_2857, n_2858, n_2859, n_2860, n_2861, n_2862, n_2863, n_2864;
  wire n_2865, n_2866, n_2867, n_2868, n_2869, n_2870, n_2871, n_2872;
  wire n_2873, n_2874, n_2875, n_2876, n_2877, n_2878, n_2879, n_2880;
  wire n_2881, n_2882, n_2883, n_2884, n_2885, n_2886, n_2887, n_2888;
  wire n_2889, n_2890, n_2891, n_2892, n_2893, n_2894, n_2895, n_2896;
  wire n_2897, n_2898, n_2899, n_2900, n_2901, n_2902, n_2903, n_2904;
  wire n_2905, n_2906, n_2907, n_2908, n_2909, n_2910, n_2911, n_2912;
  wire n_2913, n_2914, n_2915, n_2916, n_2917, n_2918, n_2919, n_2920;
  wire n_2921, n_2922, n_2923, n_2924, n_2925, n_2926, n_2927, n_2928;
  wire n_2929, n_2930, n_2931, n_2932, n_2933, n_2934, n_2935, n_2936;
  wire n_2937, n_2938, n_2939, n_2940, n_2941, n_2942, n_2943, n_2944;
  wire n_2945, n_2946, n_2947, n_2948, n_2949, n_2950, n_2951, n_2952;
  wire n_2953, n_2954, n_2955, n_2956, n_2957, n_2958, n_2959, n_2960;
  wire n_2961, n_2962, n_2963, n_2964, n_2965, n_2966, n_2967, n_2968;
  wire n_2969, n_2970, n_2971, n_2972, n_2973, n_2974, n_2975, n_2976;
  wire n_2977, n_2978, n_2979, n_2980, n_2981, n_2982, n_2983, n_2984;
  wire n_2985, n_2986, n_2987, n_2988, n_2989, n_2990, n_2991, n_2992;
  wire n_2993, n_2995, n_2996, n_2997, n_2998, n_2999, n_3000, n_3001;
  wire n_3002, n_3003, n_3004, n_3005, n_3006, n_3007, n_3008, n_3009;
  wire n_3010, n_3011, n_3012, n_3013, n_3014, n_3015, n_3016, n_3017;
  wire n_3018, n_3019, n_3020, n_3021, n_3022, n_3023, n_3024, n_3025;
  wire n_3026, n_3027, n_3028, n_3029, n_3030, n_3031, n_3032, n_3033;
  wire n_3034, n_3035, n_3036, n_3037, n_3038, n_3039, n_3040, n_3041;
  wire n_3043, n_3044, n_3045, n_3046, n_3047, n_3048, n_3049, n_3050;
  wire n_3051, n_3052, n_3053, n_3054, n_3055, n_3056, n_3057, n_3058;
  wire n_3059, n_3065, n_3066, n_3067, n_3068, n_3069, n_3070, n_3071;
  wire n_3072, n_3073, n_3074, n_3075, n_3076, n_3077, n_3078, n_3079;
  wire n_3080, n_3081, n_3082, n_3083, n_3084, n_3085, n_3086, n_3087;
  wire n_3088, n_3089, n_3090, n_3091, n_3092, n_3093, n_3094, n_3095;
  wire n_3096, n_3097, n_3098, n_3099, n_3100, n_3101, n_3102, n_3103;
  wire n_3104, n_3105, n_3106, n_3107, n_3108, n_3109, n_3110, n_3111;
  wire n_3112, n_3113, n_3114, n_3115, n_3116, n_3117, n_3118, n_3119;
  wire n_3120, n_3121, n_3122, n_3123, n_3124, n_3125, n_3126, n_3127;
  wire n_3128, n_3129, n_3130, n_3131, n_3132, n_3133, n_3134, n_3135;
  wire n_3136, n_3137, n_3138, n_3139, n_3140, n_3141, n_3142, n_3143;
  wire n_3144, n_3145, n_3146, n_3147, n_3148, n_3149, n_3150, n_3151;
  wire n_3152, n_3153, n_3154, n_3155, n_3156, n_3157, n_3158, n_3159;
  wire n_3160, n_3161, n_3162, n_3163, n_3164, n_3165, n_3166, n_3167;
  wire n_3168, n_3169, n_3170, n_3171, n_3172, n_3173, n_3174, n_3175;
  wire n_3176, n_3177, n_3178, n_3179, n_3180, n_3181, n_3182, n_3183;
  wire n_3184, n_3185, n_3186, n_3187, n_3188, n_3189, n_3190, n_3191;
  wire n_3192, n_3193, n_3194, n_3195, n_3196, n_3197, n_3198, n_3199;
  wire n_3200, n_3201, n_3202, n_3203, n_3204, n_3205, n_3206, n_3207;
  wire n_3208, n_3209, n_3210, n_3212, n_3213, n_3214, n_3215, n_3216;
  wire n_3217, n_3218, n_3219, n_3220, n_3221, n_3225, n_3226, n_3229;
  wire n_3233, n_3236, n_3237, n_3238, n_3239, n_3240, n_3241, n_3242;
  wire n_3243, n_3244, n_3245, n_3246, n_3247, n_3248, n_3249, n_3250;
  wire n_3251, n_3252, n_3253, n_3254, n_3255, n_3256, n_3257, n_3258;
  wire n_3259, n_3260, n_3261, n_3262, n_3263, n_3264, n_3265, n_3266;
  wire n_3267, n_3268, n_3269, n_3270, n_3271, n_3272, n_3273, n_3274;
  wire n_3275, n_3276, n_3277, n_3278, n_3279, n_3280, n_3281, n_3282;
  wire n_3283, n_3284, n_3285, n_3286, n_3287, n_3288, n_3289, n_3290;
  wire n_3291, n_3292, n_3293, n_3294, n_3295, n_3296, n_3297, n_3298;
  wire n_3299, n_3300, n_3301, n_3302, n_3303, n_3304, n_3305, n_3306;
  wire n_3307, n_3308, n_3309, n_3310, n_3311, n_3312, n_3313, n_3314;
  wire n_3315, n_3316, n_3317, n_3318, n_3319, n_3320, n_3321, n_3322;
  wire n_3323, n_3324, n_3325, n_3326, n_3327, n_3328, n_3329, n_3330;
  wire n_3331, n_3332, n_3333, n_3334, n_3335, n_3336, n_3337, n_3338;
  wire n_3339, n_3340, n_3341, n_3342, n_3343, n_3344, n_3345, n_3346;
  wire n_3347, n_3348, n_3349, n_3350, n_3351, n_3352, n_3353, n_3354;
  wire n_3355, n_3356, n_3357, n_3358, n_3359, n_3360, n_3361, n_3362;
  wire n_3363, n_3364, n_3365, n_3366, n_3367, n_3368, n_3369, n_3370;
  wire n_3371, n_3372, n_3373, n_3374, n_3375, n_3376, n_3377, n_3378;
  wire n_3379, n_3380, n_3381, n_3382, n_3383, n_3384, n_3385, n_3386;
  wire n_3387, n_3388, n_3389, n_3390, n_3391, n_3392, n_3393, n_3394;
  wire n_3395, n_3396, n_3397, n_3398, n_3399, n_3400, n_3401, n_3402;
  wire n_3403, n_3404, n_3405, n_3406, n_3407, n_3408, n_3409, n_3410;
  wire n_3411, n_3412, n_3413, n_3414, n_3415, n_3416, n_3417, n_3418;
  wire n_3419, n_3420, n_3421, n_3422, n_3423, n_3424, n_3425, n_3426;
  wire n_3427, n_3428, n_3429, n_3430, n_3431, n_3432, n_3433, n_3465;
  wire n_3466, n_3467, n_3468, n_3469, n_3470, n_3471, n_3472, n_3473;
  wire n_3474, n_3475, n_3476, n_3477, n_3478, n_3479, n_3480, n_3481;
  wire n_3482, n_3483, n_3484, n_3485, n_3486, n_3487, n_3488, n_3489;
  wire n_3490, n_3491, n_3492, n_3493, n_3494, n_3495, n_3496, n_3497;
  wire n_3498, n_3499, n_3500, n_3501, n_3502, n_3503, n_3504, n_3505;
  wire n_3506, n_3507, n_3508, n_3509, n_3510, n_3511, n_3512, n_3513;
  wire n_3514, n_3515, n_3516, n_3517, n_3518, n_3519, n_3520, n_3521;
  wire n_3522, n_3523, n_3524, n_3525, n_3526, n_3527, n_3528, n_3529;
  wire n_3530, n_3531, n_3532, n_3533, n_3534, n_3535, n_3536, n_3537;
  wire n_3538, n_3539, n_3540, n_3541, n_3542, n_3543, n_3544, n_3545;
  wire n_3546, n_3547, n_3548, n_3549, n_3550, n_3551, n_3552, n_3553;
  wire n_3554, n_3555, n_3556, n_3557, n_3558, n_3559, n_3560, n_3561;
  wire n_3562, n_3563, n_3564, n_3565, n_3566, n_3567, n_3568, n_3569;
  wire n_3570, n_3571, n_3572, n_3573, n_3574, n_3575, n_3576, n_3577;
  wire n_3578, n_3579, n_3580, n_3581, n_3582, n_3583, n_3584, n_3585;
  wire n_3586, n_3587, n_3588, n_3589, n_3590, n_3591, n_3592, n_3593;
  wire n_3594, n_3595, n_3596, n_3597, n_3598, n_3599, n_3600, n_3601;
  wire n_3602, n_3603, n_3604, n_3605, n_3606, n_3607, n_3608, n_3609;
  wire n_3610, n_3611, n_3612, n_3613, n_3614, n_3615, n_3616, n_3617;
  wire n_3618, n_3619, n_3620, n_3621, n_3622, n_3623, n_3624, n_3625;
  wire n_3626, n_3627, n_3628, n_3629, n_3630, n_3631, n_3632, n_3633;
  wire n_3634, n_3635, n_3636, n_3637, n_3638, n_3639, n_3640, n_3641;
  wire n_3642, n_3643, n_3644, n_3645, n_3646, n_3647, n_3648, n_3649;
  wire n_3650, n_3651, n_3652, n_3653, n_3654, n_3655, n_3656, n_3657;
  wire n_3658, n_3659, n_3660, n_3661, n_3662, n_3663, n_3664, n_3665;
  wire n_3666, n_3667, n_3668, n_3669, n_3670, n_3671, n_3672, n_3673;
  wire n_3674, n_3675, n_3676, n_3677, n_3678, n_3679, n_3680, n_3681;
  wire n_3682, n_3683, n_3684, n_3685, n_3686, n_3687, n_3688, n_3689;
  wire n_3690, n_3691, n_3692, n_3693, n_3694, n_3695, n_3696, n_3697;
  wire n_3698, n_3699, n_3700, n_3701, n_3702, n_3703, n_3704, n_3705;
  wire n_3706, n_3707, n_3708, n_3709, n_3710, n_3711, n_3712, n_3713;
  wire n_3714, n_3715, n_3716, n_3717, n_3718, n_3719, n_3720, n_3721;
  wire n_3722, n_3723, n_3724, n_3725, n_3726, n_3727, n_3728, n_3729;
  wire n_3730, n_3731, n_3732, n_3733, n_3734, n_3735, n_3736, n_3737;
  wire n_3738, n_3739, n_3740, n_3741, n_3742, n_3743, n_3744, n_3745;
  wire n_3746, n_3747, n_3748, n_3749, n_3750, n_3751, n_3752, n_3753;
  wire n_3754, n_3755, n_3756, n_3757, n_3758, n_3759, n_3760, n_3761;
  wire n_3762, n_3763, n_3764, n_3765, n_3766, n_3767, n_3768, n_3769;
  wire n_3770, n_3771, n_3772, n_3773, n_3774, n_3775, n_3776, n_3777;
  wire n_3778, n_3779, n_3780, n_3781, n_3782, n_3783, n_3784, n_3785;
  wire n_3786, n_3787, n_3788, n_3789, n_3790, n_3791, n_3792, n_3793;
  wire n_3794, n_3795, n_3796, n_3797, n_3798, n_3799, n_3800, n_3801;
  wire n_3802, n_3803, n_3804, n_3805, n_3806, n_3807, n_3808, n_3809;
  wire n_3810, n_3811, n_3812, n_3813, n_3814, n_3815, n_3816, n_3817;
  wire n_3818, n_3819, n_3820, n_3821, n_3822, n_3823, n_3824, n_3825;
  wire n_3826, n_3827, n_3828, n_3829, n_3830, n_3831, n_3832, n_3833;
  wire n_3834, n_3835, n_3836, n_3837, n_3838, n_3839, n_3840, n_3841;
  wire n_3842, n_3843, n_3844, n_3845, n_3846, n_3847, n_3848, n_3849;
  wire n_3850, n_3851, n_3852, n_3853, n_3854, n_3855, n_3856, n_3857;
  wire n_3858, n_3859, n_3860, n_3861, n_3862, n_3863, n_3864, n_3865;
  wire n_3866, n_3867, n_3868, n_3869, n_3870, n_3871, n_3872, n_3873;
  wire n_3874, n_3875, n_3876, n_3877, n_3878, n_3879, n_3880, n_3881;
  wire n_3882, n_3883, n_3884, n_3885, n_3886, n_3887, n_3888, n_3889;
  wire n_3890, n_3891, n_3892, n_3893, n_3894, n_3895, n_3896, n_3897;
  wire n_3898, n_3899, n_3900, n_3901, n_3902, n_3903, n_3904, n_3905;
  wire n_3906, n_3907, n_3908, n_3909, n_3910, n_3911, n_3912, n_3913;
  wire n_3914, n_3915, n_3916, n_3917, n_3918, n_3919, n_3920, n_3921;
  wire n_3922, n_3923, n_3924, n_3925, n_3926, n_3927, n_3928, n_3929;
  wire n_3930, n_3931, n_3932, n_3933, n_3934, n_3935, n_3936, n_3937;
  wire n_3938, n_3939, n_3940, n_3941, n_3942, n_3943, n_3944, n_3945;
  wire n_3946, n_3947, n_3948, n_3949, n_3950, n_3951, n_3952, n_3953;
  wire n_3954, n_3955, n_3956, n_3957, n_3958, n_3959, n_3960, n_3961;
  wire n_3962, n_3963, n_3964, n_3965, n_3966, n_3967, n_3968, n_3969;
  wire n_3970, n_3971, n_3972, n_3973, n_3974, n_3975, n_3976, n_3977;
  wire n_3978, n_3979, n_3980, n_3981, n_3982, n_3983, n_3984, n_3985;
  wire n_3986, n_3987, n_3988, n_3989, n_3990, n_3991, n_3992, n_3993;
  wire n_3994, n_3995, n_3996, n_3997, n_3998, n_3999, n_4000, n_4001;
  wire n_4002, n_4003, n_4004, n_4005, n_4006, n_4007, n_4008, n_4009;
  wire n_4010, n_4011, n_4012, n_4013, n_4014, n_4015, n_4016, n_4017;
  wire n_4018, n_4019, n_4020, n_4021, n_4022, n_4023, n_4024, n_4025;
  wire n_4026, n_4027, n_4028, n_4029, n_4030, n_4031, n_4032, n_4033;
  wire n_4034, n_4035, n_4036, n_4037, n_4038, n_4039, n_4040, n_4041;
  wire n_4042, n_4043, n_4044, n_4045, n_4046, n_4047, n_4048, n_4049;
  wire n_4050, n_4051, n_4052, n_4053, n_4054, n_4055, n_4056, n_4057;
  wire n_4058, n_4059, n_4060, n_4061, n_4062, n_4063, n_4064, n_4065;
  wire n_4066, n_4067, n_4068, n_4069, n_4070, n_4071, n_4072, n_4073;
  wire n_4074, n_4075, n_4076, n_4077, n_4078, n_4079, n_4080, n_4081;
  wire n_4082, n_4083, n_4084, n_4085, n_4086, n_4087, n_4088, n_4089;
  wire n_4090, n_4091, n_4092, n_4093, n_4094, n_4095, n_4096, n_4097;
  wire n_4098, n_4099, n_4100, n_4101, n_4102, n_4103, n_4104, n_4105;
  wire n_4106, n_4107, n_4108, n_4109, n_4110, n_4111, n_4112, n_4113;
  wire n_4114, n_4115, n_4116, n_4117, n_4118, n_4119, n_4120, n_4121;
  wire n_4122, n_4123, n_4124, n_4125, n_4126, n_4127, n_4128, n_4129;
  wire n_4130, n_4131, n_4132, n_4133, n_4134, n_4135, n_4136, n_4137;
  wire n_4138, n_4139, n_4140, n_4141, n_4142, n_4143, n_4144, n_4145;
  wire n_4146, n_4147, n_4148, n_4149, n_4150, n_4151, n_4152, n_4153;
  wire n_4154, n_4155, n_4156, n_4157, n_4158, n_4159, n_4160, n_4161;
  wire n_4162, n_4163, n_4164, n_4165, n_4166, n_4167, n_4168, n_4169;
  wire n_4170, n_4171, n_4172, n_4173, n_4174, n_4175, n_4176, n_4177;
  wire n_4178, n_4179, n_4180, n_4181, n_4182, n_4183, n_4184, n_4185;
  wire n_4186, n_4187, n_4188, n_4189, n_4190, n_4191, n_4192, n_4193;
  wire n_4194, n_4195, n_4196, n_4197, n_4198, n_4199, n_4200, n_4201;
  wire n_4202, n_4203, n_4204, n_4205, n_4206, n_4207, n_4208, n_4209;
  wire n_4210, n_4211, n_4212, n_4213, n_4214, n_4215, n_4216, n_4217;
  wire n_4218, n_4219, n_4220, n_4221, n_4222, n_4223, n_4224, n_4225;
  wire n_4226, n_4227, n_4228, n_4229, n_4230, n_4231, n_4232, n_4233;
  wire n_4234, n_4235, n_4236, n_4237, n_4238, n_4239, n_4240, n_4241;
  wire n_4242, n_4243, n_4244, n_4245, n_4246, n_4247, n_4248, n_4249;
  wire n_4250, n_4251, n_4252, n_4253, n_4254, n_4255, n_4256, n_4257;
  wire n_4258, n_4259, n_4260, n_4261, n_4262, n_4263, n_4264, n_4265;
  wire n_4266, n_4267, n_4268, n_4269, n_4270, n_4271, n_4272, n_4273;
  wire n_4274, n_4275, n_4276, n_4277, n_4278, n_4279, n_4280, n_4281;
  wire n_4282, n_4287, n_4288, n_4289, n_4290, n_4291, n_4292, n_4293;
  wire n_4294, n_4295, n_4296, n_4297, n_4298, n_4299, n_4300, n_4301;
  wire n_4302, n_4303, n_4304, n_4305, n_4306, n_4307, n_4308, n_4309;
  wire n_4310, n_4311, n_4312, n_4313, n_4314, n_4315, n_4316, n_4317;
  wire n_4318, n_4319, n_4320, n_4321, n_4322, n_4323, n_4324, n_4325;
  wire n_4326, n_4327, n_4328, n_4329, n_4330, n_4331, n_4332, n_4333;
  wire n_4334, n_4335, n_4336, n_4337, n_4338, n_4339, n_4340, n_4341;
  wire n_4342, n_4343, n_4344, n_4345, n_4346, n_4347, n_4348, n_4349;
  wire n_4350, n_4351, n_4352, n_4353, n_4354, n_4355, n_4356, n_4357;
  wire n_4358, n_4359, n_4360, n_4361, n_4362, n_4363, n_4364, n_4365;
  wire n_4366, n_4367, n_4368, n_4369, n_4370, n_4371, n_4372, n_4373;
  wire n_4374, n_4375, n_4376, n_4377, n_4378, n_4379, n_4380, n_4381;
  wire n_4382, n_4383, n_4384, n_4385, n_4386, n_4387, n_4388, n_4389;
  wire n_4390, n_4391, n_4392, n_4393, n_4394, n_4395, n_4396, n_4397;
  wire n_4398, n_4399, n_4400, n_4401, n_4402, n_4403, n_4404, n_4405;
  wire n_4406, n_4407, n_4408, n_4409, n_4410, n_4411, n_4412, n_4413;
  wire n_4414, n_4415, n_4416, n_4417, n_4418, n_4419, n_4420, n_4421;
  wire n_4422, n_4423, n_4424, n_4425, n_4426, n_4427, n_4428, n_4429;
  wire n_4430, n_4431, n_4432, n_4433, n_4434, n_4435, n_4436, n_4437;
  wire n_4438, n_4439, n_4440, n_4441, n_4442, n_4443, n_4444, n_4445;
  wire n_4446, n_4447, n_4448, n_4449, n_4450, n_4451, n_4452, n_4453;
  wire n_4454, n_4455, n_4456, n_4457, n_4458, n_4459, n_4460, n_4461;
  wire n_4462, n_4463, n_4464, n_4465, n_4466, n_4467, n_4468, n_4469;
  wire n_4470, n_4471, n_4472, n_4473, n_4474, n_4475, n_4476, n_4477;
  wire n_4478, n_4479, n_4480, n_4481, n_4482, n_4483, n_4484, n_4485;
  wire n_4486, n_4487, n_4488, n_4489, n_4490, n_4491, n_4492, n_4493;
  wire n_4494, n_4495, n_4496, n_4497, n_4498, n_4499, n_4500, n_4501;
  wire n_4502, n_4503, n_4504, n_4505, n_4506, n_4507, n_4508, n_4509;
  wire n_4510, n_4511, n_4512, n_4513, n_4514, n_4515, n_4516, n_4517;
  wire n_4518, n_4519, n_4520, n_4521, n_4522, n_4523, n_4524, n_4525;
  wire n_4526, n_4527, n_4528, n_4529, n_4530, n_4531, n_4532, n_4533;
  wire n_4534, n_4535, n_4536, n_4537, n_4538, n_4539, n_4540, n_4541;
  wire n_4542, n_4543, n_4544, n_4545, n_4546, n_4547, n_4548, n_4549;
  wire n_4550, n_4551, n_4552, n_4553, n_4554, n_4555, n_4556, n_4557;
  wire n_4558, n_4559, n_4560, n_4561, n_4562, n_4563, n_4564, n_4565;
  wire n_4566, n_4567, n_4568, n_4569, n_4570, n_4571, n_4572, n_4573;
  wire n_4574, n_4575, n_4576, n_4577, n_4578, n_4579, n_4580, n_4581;
  wire n_4582, n_4583, n_4584, n_4585, n_4586, n_4587, n_4588, n_4589;
  wire n_4590, n_4591, n_4592, n_4593, n_4594, n_4595, n_4596, n_4597;
  wire n_4598, n_4599, n_4600, n_4601, n_4602, n_4603, n_4604, n_4605;
  wire n_4606, n_4607, n_4608, n_4609, n_4610, n_4611, n_4612, n_4613;
  wire n_4614, n_4615, n_4616, n_4617, n_4618, n_4619, n_4620, n_4621;
  wire n_4622, n_4623, n_4624, n_4625, n_4626, n_4627, n_4628, n_4629;
  wire n_4630, n_4631, n_4632, n_4633, n_4634, n_4635, n_4636, n_4637;
  wire n_4638, n_4639, n_4640, n_4641, n_4642, n_4643, n_4644, n_4645;
  wire n_4646, n_4647, n_4648, n_4649, n_4650, n_4651, n_4652, n_4653;
  wire n_4654, n_4655, n_4656, n_4657, n_4658, n_4659, n_4660, n_4661;
  wire n_4662, n_4663, n_4664, n_4665, n_4666, n_4667, n_4668, n_4669;
  wire n_4670, n_4671, n_4672, n_4673, n_4674, n_4675, n_4676, n_4677;
  wire n_4678, n_4679, n_4680, n_4681, n_4682, n_4683, n_4684, n_4685;
  wire n_4686, n_4687, n_4688, n_4689, n_4690, n_4691, n_4692, n_4693;
  wire n_4694, n_4695, n_4696, n_4697, n_4698, n_4699, n_4700, n_4701;
  wire n_4702, n_4703, n_4704, n_4705, n_4706, n_4707, n_4708, n_4709;
  wire n_4710, n_4712, n_4713, n_4714, n_4715, n_4716, n_4717, n_4718;
  wire n_4719, n_4720, n_4721, n_4722, n_4723, n_4724, n_4725, n_4726;
  wire n_4727, n_4728, n_4729, n_4730, n_4731, n_4732, n_4733, n_4734;
  wire n_4735, n_4736, n_4737, n_4738, n_4739, n_4740, n_4741, n_4742;
  wire n_4743, n_4744, n_4745, n_4746, n_4747, n_4748, n_4749, n_4750;
  wire n_4751, n_4752, n_4753, n_4754, n_4755, n_4756, n_4757, n_4758;
  wire n_4759, n_4760, n_4761, n_4762, n_4763, n_4764, n_4765, n_4766;
  wire n_4767, n_4768, n_4769, n_4770, n_4771, n_4772, n_4773, n_4774;
  wire n_4775, n_4776, n_4777, n_4778, n_4779, n_4780, n_4781, n_4782;
  wire n_4783, n_4784, n_4785, n_4786, n_4787, n_4788, n_4789, n_4790;
  wire n_4791, n_4792, n_4793, n_4794, n_4795, n_4796, n_4797, n_4798;
  wire n_4799, n_4800, n_4801, n_4802, n_4803, n_4804, n_4805, n_4806;
  wire n_4807, n_4808, n_4809, n_4810, n_4811, n_4812, n_4813, n_4814;
  wire n_4815, n_4816, n_4817, n_4818, n_4819, n_4820, n_4821, n_4822;
  wire n_4823, n_4824, n_4825, n_4826, n_4827, n_4828, n_4829, n_4830;
  wire n_4831, n_4832, n_4833, n_4834, n_4835, n_4836, n_4837, n_4838;
  wire n_4839, n_4840, n_4841, n_4842, n_4844, n_4845, n_4846, n_4847;
  wire n_4848, n_4849, n_4850, n_4851, n_4852, n_4853, n_4854, n_4855;
  wire n_4856, n_4857, n_4858, n_4859, n_4860, n_4861, n_4862, n_4863;
  wire n_4864, n_4865, n_4866, n_4867, n_4868, n_4869, n_4870, n_4871;
  wire n_4872, n_4873, n_4874, n_4875, n_4877, n_4878, n_4879, n_4880;
  wire n_4881, n_4882, n_4883, n_4884, n_4885, n_4886, n_4887, n_4888;
  wire n_4889, n_4890, n_4891, n_4892, n_4893, n_4894, n_4895, n_4896;
  wire n_4897, n_4898, n_4899, n_4900, n_4901, n_4902, n_4905, n_4906;
  wire n_4907, n_4908, n_4909, n_4910, n_4911, n_4912, n_4913, n_4914;
  wire n_4915, n_4916, n_4917, n_4918, n_4919, n_4920, n_4921, n_4922;
  wire n_4923, n_4924, n_4925, n_4926, n_4927, n_4928, n_4929, n_4930;
  wire n_4931, n_4932, n_4933, n_4934, n_4935, n_4936, n_4937, n_4938;
  wire n_4939, n_4940, n_4941, n_4942, n_4943, n_4944, n_4945, n_4946;
  wire n_4947, n_4948, n_4949, n_4950, n_4951, n_4952, n_4953, n_4954;
  wire n_4955, n_4956, n_4957, n_4958, n_4959, n_4960, n_4961, n_4962;
  wire n_4963, n_4964, n_4965, n_4966, n_4967, n_4968, n_4969, n_4970;
  wire n_4971, n_4972, n_4973, n_4974, n_4975, n_4976, n_4977, n_4978;
  wire n_4979, n_4980, n_4981, n_4982, n_4983, n_4984, n_4985, n_4986;
  wire n_4987, n_4989, n_4990, n_4991, n_4992, n_4993, n_4994, n_4995;
  wire n_4996, n_4997, n_4998, n_4999, n_5000, n_5001, n_5002, n_5003;
  wire n_5004, n_5005, n_5006, n_5007, n_5008, n_5009, n_5010, n_5011;
  wire n_5012, n_5013, n_5014, n_5015, n_5016, n_5017, n_5018, n_5019;
  wire n_5020, n_5021, n_5022, n_5023, n_5024, n_5025, n_5026, n_5027;
  wire n_5028, n_5029, n_5030, n_5031, n_5032, n_5033, n_5034, n_5035;
  wire n_5036, n_5037, n_5038, n_5039, n_5040, n_5041, n_5042, n_5043;
  wire n_5044, n_5045, n_5046, n_5047, n_5048, n_5049, n_5050, n_5051;
  wire n_5052, n_5053, n_5054, n_5055, n_5056, n_5057, n_5059, n_5060;
  wire n_5061, n_5062, n_5063, n_5064, n_5065, n_5066, n_5067, n_5068;
  wire n_5069, n_5070, n_5071, n_5072, n_5073, n_5074, n_5075, n_5076;
  wire n_5077, n_5078, n_5079, n_5080, n_5081, n_5082, n_5083, n_5084;
  wire n_5085, n_5086, n_5087, n_5088, n_5089, n_5090, n_5091, n_5092;
  wire n_5093, n_5094, n_5095, n_5096, n_5097, n_5098, n_5099, n_5100;
  wire n_5101, n_5102, n_5103, n_5104, n_5105, n_5106, n_5107, n_5108;
  wire n_5109, n_5110, n_5111, n_5112, n_5113, n_5114, n_5115, n_5116;
  wire n_5117, n_5118, n_5119, n_5120, n_5121, n_5122, n_5123, n_5124;
  wire n_5125, n_5126, n_5127, n_5128, n_5129, n_5130, n_5131, n_5132;
  wire n_5133, n_5134, n_5135, n_5136, n_5137, n_5138, n_5139, n_5140;
  wire n_5141, n_5142, n_5143, n_5144, n_5145, n_5146, n_5147, n_5148;
  wire n_5149, n_5150, n_5151, n_5152, n_5153, n_5154, n_5155, n_5156;
  wire n_5157, n_5158, n_5159, n_5160, n_5161, n_5162, n_5163, n_5164;
  wire n_5165, n_5166, n_5167, n_5168, n_5169, n_5170, n_5171, n_5172;
  wire n_5173, n_5174, n_5175, n_5176, n_5177, n_5178, n_5179, n_5180;
  wire n_5181, n_5182, n_5183, n_5184, n_5185, n_5186, n_5187, n_5188;
  wire n_5189, n_5190, n_5191, n_5192, n_5193, n_5194, n_5195, n_5196;
  wire n_5197, n_5198, n_5199, n_5200, n_5201, n_5202, n_5203, n_5204;
  wire n_5205, n_5206, n_5207, n_5208, n_5209, n_5210, n_5211, n_5212;
  wire n_5213, n_5214, n_5215, n_5216, n_5217, n_5218, n_5219, n_5220;
  wire n_5221, n_5222, n_5223, n_5224, n_5225, n_5226, n_5227, n_5228;
  wire n_5229, n_5230, n_5231, n_5232, n_5233, n_5234, n_5235, n_5236;
  wire n_5237, n_5238, n_5239, n_5240, n_5241, n_5242, n_5243, n_5244;
  wire n_5245, n_5246, n_5247, n_5248, n_5249, n_5250, n_5251, n_5252;
  wire n_5253, n_5254, n_5255, n_5256, n_5257, n_5259, n_5260, n_5261;
  wire n_5262, n_5263, n_5264, n_5265, n_5266, n_5267, n_5268, n_5269;
  wire n_5270, n_5272, n_5273, n_5274, n_5275, n_5276, n_5277, n_5278;
  wire n_5279, n_5280, n_5281, n_5282, n_5283, n_5284, n_5285, n_5286;
  wire n_5287, n_5288, n_5289, n_5290, n_5291, n_5292, n_5293, n_5294;
  wire n_5295, n_5296, n_5297, n_5298, n_5299, n_5300, n_5301, n_5302;
  wire n_5303, n_5304, n_5305, n_5306, n_5307, n_5308, n_5309, n_5310;
  wire n_5311, n_5312, n_5313, n_5314, n_5315, n_5316, n_5317, n_5318;
  wire n_5319, n_5320, n_5321, n_5322, n_5323, n_5324, n_5325, n_5326;
  wire n_5327, n_5328, n_5329, n_5330, n_5331, n_5332, n_5333, n_5334;
  wire n_5335, n_5336, n_5337, n_5338, n_5339, n_5340, n_5341, n_5342;
  wire n_5343, n_5344, n_5345, n_5346, n_5347, n_5348, n_5349, n_5350;
  wire n_5351, n_5352, n_5353, n_5354, n_5355, n_5356, n_5357, n_5358;
  wire n_5359, n_5360, n_5361, n_5362, n_5363, n_5364, n_5365, n_5366;
  wire n_5398, n_5399, n_5400, n_5401, n_5402, n_5403, n_5404, n_5405;
  wire n_5406, n_5407, n_5408, n_5409, n_5410, n_5411, n_5412, n_5413;
  wire n_5414, n_5415, n_5416, n_5417, n_5418, n_5419, n_5420, n_5421;
  wire n_5422, n_5423, n_5424, n_5425, n_5426, n_5427, n_5428, n_5429;
  wire n_5431, n_5432, n_5433, n_5434, n_5435, n_5436, n_5437, n_5438;
  wire n_5439, n_5440, n_5441, n_5442, n_5443, n_5444, n_5445, n_5446;
  wire n_5447, n_5448, n_5449, n_5450, n_5451, n_5452, n_5453, n_5454;
  wire n_5455, n_5456, n_5457, n_5458, n_5459, n_5460, n_5461, n_5462;
  wire n_5463, n_5464, n_5465, n_5466, n_5467, n_5468, n_5469, n_5470;
  wire n_5471, n_5472, n_5473, n_5474, n_5475, n_5476, n_5477, n_5478;
  wire n_5479, n_5480, n_5481, n_5482, n_5483, n_5484, n_5485, n_5486;
  wire n_5487, n_5488, n_5489, n_5490, n_5491, n_5492, n_5493, n_5494;
  wire n_5495, n_5496, n_5497, n_5498, n_5499, n_5500, n_5501, n_5502;
  wire n_5503, n_5504, n_5505, n_5506, n_5507, n_5508, n_5509, n_5510;
  wire n_5511, n_5512, n_5513, n_5514, n_5515, n_5516, n_5517, n_5518;
  wire n_5519, n_5520, n_5521, n_5522, n_5523, n_5524, n_5525, n_5526;
  wire n_5527, n_5528, n_5585, n_5586, n_5587, n_5588, n_5589, n_5590;
  wire n_5591, n_5592, n_5593, n_5594, n_5595, n_5596, n_5597, n_5598;
  wire n_5599, n_5600, n_5601, n_5602, n_5603, n_5604, n_5605, n_5606;
  wire n_5607, n_5608, n_5609, n_5610, n_5611, n_5612, n_5613, n_5614;
  wire n_5615, n_5616, n_5617, n_5626, n_5627, n_5628, n_5629, n_5630;
  wire n_5631, n_5632, n_5633, n_5634, n_5635, n_5636, n_5637, n_5638;
  wire n_5639, n_5640, n_5641, n_5642, n_5643, n_5644, n_5645, n_5646;
  wire n_5647, n_5648, n_5649, n_5650, n_5651, n_5652, n_5653, n_5654;
  wire n_5655, n_5656, n_5657, n_5658, n_5659, n_5660, n_5661, n_5662;
  wire n_5663, n_5664, n_5665, n_5666, n_5667, n_5668, n_5669, n_5670;
  wire n_5671, n_5672, n_5673, n_5674, n_5675, n_5676, n_5677, n_5678;
  wire n_5679, n_5680, n_5681, n_5682, n_5683, n_5684, n_5685, n_5686;
  wire n_5687, n_5688, n_5689, n_5690, n_5691, n_5692, n_5693, n_5694;
  wire n_5784, n_5786, n_5788, n_5813, n_5827, n_5829, n_5859, n_5970;
  wire n_5974, n_5980, n_5984, n_5993, n_5994, n_5995, n_5996, n_5997;
  wire n_5998, n_5999, n_6011, n_6026, n_6027, n_6028, n_6029, n_6030;
  wire n_6031, n_6032, n_6033, n_6034, n_6035, n_6036, n_6037, n_6038;
  wire n_6039, n_6040, n_6041, n_6042, n_6043, n_6044, n_6045, n_6048;
  wire n_6050, n_6051, n_6052, n_6053, n_6054, n_6055, n_6056, n_6057;
  wire n_6058, n_6059, n_6060, n_6061, n_6063, n_6064, n_6066, n_6067;
  wire n_6068, n_6070, n_6071, n_6072, n_6073, n_6082, n_6083, n_6084;
  wire n_6085, n_6086, n_6087, n_6088, n_6089, n_6090, n_6091, n_6092;
  wire n_6093, n_6094, n_6095, n_6096, n_6097, n_6098, n_6099, n_6100;
  wire n_6101, n_6102, n_6103, n_6104, n_6105, n_6106, n_6110, n_6111;
  wire n_6112, n_6113, n_6114, n_6115, n_6117, n_6118, n_6119, n_6121;
  wire n_6122, n_6124, n_6127, n_6128, n_6129, n_6130, n_6131, n_6132;
  wire n_6133, n_6134, n_6135, n_6136, n_6137, n_6138, n_6140, n_6141;
  wire n_6142, n_6143, n_6144, n_6145, n_6146, n_6147, n_6148, n_6149;
  wire n_6150, n_6151, n_6152, n_6160, n_6161, n_6162, n_6165, n_6166;
  wire n_6167, n_6168, n_6169, n_6170, n_6171, n_6172, n_6173, n_6175;
  wire n_6176, n_6177, n_6178, n_6179, n_6181, n_6182, n_6183, n_6184;
  wire n_6185, n_6186, n_6187, n_6188, n_6189, n_6190, n_6191, n_6192;
  wire n_6193, n_6195, n_6196, n_6201, n_6208, n_6211, n_6212, n_6213;
  wire n_6214, n_6215, n_6216, n_6217, n_6218, n_6219, n_6220, n_6222;
  wire n_6223, n_6224, n_6227, n_6228, n_6229, n_6230, n_6231, n_6232;
  wire n_6233, n_6234, n_6235, n_6236, n_6237, n_6238, n_6239, n_6240;
  wire n_6241, n_6242, n_6243, n_6244, n_6245, n_6246, n_6247, n_6248;
  wire n_6249, n_6250, n_6251, n_6252, n_6253, n_6254, n_6255, n_6256;
  wire n_6257, n_6258, n_6259, n_6260, n_6266, n_6270, n_6271, n_6272;
  wire n_6273, n_6274, n_6275, n_6276, n_6278, n_6280, n_6282, n_6283;
  wire n_6284, n_6285, n_6287, n_6288, n_6289, n_6290, n_6291, n_6292;
  wire n_6293, n_6294, n_6295, n_6296, n_6297, n_6298, n_6299, n_6300;
  wire n_6301, n_6302, n_6303, n_6304, n_6307, n_6309, n_6310, n_6311;
  wire n_6312, n_6313, n_6314, n_6315, n_6316, n_6317, n_6318, n_6319;
  wire n_6320, n_6321, n_6322, n_6323, n_6324, n_6325, n_6326, n_6327;
  wire n_6328, n_6329, n_6330, n_6331, n_6332, n_6333, n_6334, n_6335;
  wire n_6336, n_6337, n_6338, n_6339, n_6340, n_6341, n_6342, n_6343;
  wire n_6344, n_6345, n_6346, n_6347, n_6348, n_6349, n_6350, n_6351;
  wire n_6352, n_6353, n_6365, n_6369, n_6371, n_6372, n_6514, n_6517;
  wire n_6524, n_6527, n_6530, n_6531, n_6532, n_6533, n_6534, n_6535;
  wire n_6536, n_6537, n_6538, n_6541, n_6542, n_6543, n_6544, n_6546;
  wire n_6547, n_6548, n_6549, n_6550, n_6551, n_6552, n_6553, n_6554;
  wire n_6555, n_6559, n_6565, n_6567, n_6574, n_6575, n_6576, n_6577;
  wire n_6578, n_6579, n_6580, n_6581, n_6582, n_6583, n_6584, n_6585;
  wire n_6586, n_6587, n_6588, n_6589, n_6590, n_6591, n_6592, n_6593;
  wire n_6594, n_6595, n_6596, n_6597, n_6598, n_6599, n_6600, n_6601;
  wire n_6602, n_6603, n_6604, n_6605, n_6606, n_6607, n_6608, n_6609;
  wire n_6610, n_6611, n_6612, n_6613, n_6614, n_6615, n_6616, n_6617;
  wire n_6618, n_6619, n_6620, n_6621, n_6622, n_6623, n_6624, n_6625;
  wire n_6626, n_6627, n_6628, n_6629, n_6630, n_6631, n_6632, n_6633;
  wire n_6634, n_6635, n_6636, n_6637, n_6638, n_6639, n_6640, n_6641;
  wire n_6642, n_6643, n_6644, n_6645, n_6646, n_6647, n_6648, n_6649;
  wire n_6650, n_6651, n_6652, n_6653, n_6654, n_6655, n_6656, n_6657;
  wire n_6658, n_6659, n_6660, n_6661, n_6663, n_6665, n_6666, n_6667;
  wire n_6668, n_6671, n_6672, n_6673, n_6674, n_6678, n_6679, n_6680;
  wire n_6681, n_6682, n_6683, n_6684, n_6685, n_6686, n_6687, n_6688;
  wire n_6689, n_6690, n_6691, n_6692, n_6693, n_6694, n_6695, n_6696;
  wire n_6697, n_6698, n_6699, n_6700, n_6701, n_6702, n_6703, n_6704;
  wire n_6705, n_6706, n_6707, n_6708, n_6740, n_6741, n_6742, n_6743;
  wire n_6744, n_6745, n_6746, n_6747, n_6748, n_6749, n_6750, n_6751;
  wire n_6752, n_6753, n_6754, n_6755, n_6756, n_6757, n_6758, n_6759;
  wire n_6760, n_6761, n_6762, n_6763, n_6764, n_6765, n_6766, n_6767;
  wire n_6768, n_6769, n_6770, n_6771, n_6772, n_6773, n_6774, n_6775;
  wire n_6776, n_6777, n_6778, n_6779, n_6780, n_6781, n_6782, n_6783;
  wire n_6784, n_6785, n_6786, n_6787, n_6788, n_6789, n_6790, n_6791;
  wire n_6792, n_6793, n_6794, n_6795, n_6796, n_6797, n_6798, n_6799;
  wire n_6800, n_6801, n_6802, n_6803, n_6804, n_6805, n_6806, n_6807;
  wire n_6808, n_6809, n_6810, n_6811, n_6812, n_6813, n_6814, n_6815;
  wire n_6816, n_6817, n_6819, n_6821, n_6824, n_6827, n_6828, n_6832;
  wire n_6833, n_6834, n_6835, n_6836, n_6837, n_6838, n_6839, n_6840;
  wire n_6841, n_6842, n_6843, n_6844, n_6845, n_6846, n_6847, n_6848;
  wire n_6849, n_6850, n_6851, n_6852, n_6853, n_6854, n_6855, n_6856;
  wire n_6857, n_6858, n_6859, n_6860, n_6861, n_6862, n_6864, n_6865;
  wire n_6931, n_6932, n_6933, n_6934, n_6935, n_6936, n_6937, n_6938;
  wire n_6939, n_6940, n_6941, n_6943, n_6944, n_6945, n_6947, n_6948;
  wire n_6949, n_6950, n_6951, n_6952, n_6953, n_6954, n_6955, n_6956;
  wire n_6960, n_6976, n_6985, n_6986, n_6987, n_6988, n_6989, n_6990;
  wire n_6992, n_6993, n_6994, n_6995, n_6996, n_6997, n_6998, n_6999;
  wire n_7000, n_7001, n_7002, n_7003, n_7004, n_7005, n_7006, n_7007;
  wire n_7008, n_7009, n_7010, n_7011, n_7012, n_7013, n_7014, n_7015;
  wire n_7016, n_7017, n_7018, n_7019, n_7020, n_7021, n_7022, n_7023;
  wire n_7024, n_7025, n_7026, n_7027, n_7028, n_7029, n_7030, n_7031;
  wire n_7032, n_7033, n_7034, n_7035, n_7036, n_7037, n_7038, n_7039;
  wire n_7040, n_7041, n_7042, n_7043, n_7044, n_7045, n_7046, n_7047;
  wire n_7048, n_7049, n_7050, n_7051, n_7052, n_7053, n_7054, n_7126;
  wire n_7130, n_7137, n_7139, n_7145, n_7146, n_7147, n_8138, n_8325;
  wire n_8490, n_8493, n_8514, n_8535, n_8553, n_8556, n_8577, n_8595;
  wire n_8598, n_8619, n_8640, n_8658, n_8661, n_8682, n_8703, n_8721;
  wire n_8724, n_8745, n_8766, n_8784, n_8787, n_8808, n_8829, n_8847;
  wire n_8850, n_8868, n_8871, n_8892, n_8910, n_8913, n_8931, n_8934;
  wire n_8952, n_8955, n_8976, n_8994, n_8997, n_9018, n_9039, n_9060;
  wire n_9078, n_9081, n_9099, n_9102, n_9120, n_9123, n_9141, n_9144;
  wire n_9162, n_9165, n_9183, n_9186, n_9204, n_9207, n_9225, n_9228;
  wire n_9246, n_9249, n_9267, n_9270, n_9288, n_9291, n_9309, n_9312;
  wire n_9330, n_9333, n_9351, n_9354, n_9372, n_9375, n_9393, n_9396;
  wire n_9414, n_9417, n_9435, n_9438, n_9456, n_9459, n_9477, n_9480;
  wire n_9498, n_9501, n_9519, n_9522, n_9540, n_9543, n_9564, n_9585;
  wire n_9606, n_9627, n_9648, n_9669, n_9687, n_9690, n_10451, n_10491;
  wire n_10531, n_10551, n_11689, n_11690, n_11691, n_11692, n_11693,
       n_11694;
  wire n_11695, n_11696, n_11697, n_11698, n_11699, n_11700, n_11701,
       n_11702;
  wire n_11703, n_11704, n_11705, n_11706, n_11707, n_11708, n_11709,
       n_11710;
  wire n_11711, n_11712, n_11713, n_11714, n_11715, n_11716, n_11717,
       n_11718;
  wire n_11719, n_11720, n_11721, n_11722, n_11723, n_11724, n_11725,
       n_11726;
  wire n_11727, n_11728, n_11729, n_11730, n_11731, n_11732, n_11733,
       n_11734;
  wire n_11735, n_11736, n_11737, n_11738, n_11739, n_11740, n_11741,
       n_11742;
  wire n_11743, n_11744, n_11745, n_11746, n_11747, n_11748, n_11749,
       n_11750;
  wire n_11751, n_11752, n_11753, n_11754, n_11755, n_11756, n_11757,
       n_11758;
  wire n_11759, n_11760, n_11761, n_11762, n_11763, n_11764, n_11765,
       n_11766;
  wire n_11767, n_11768, n_11769, n_11770, n_11771, n_11772, n_11773,
       n_11774;
  wire n_11775, n_11776, n_11777, n_11778, n_11779, n_11780, n_11781,
       n_11782;
  wire n_11783, n_11784, n_11785, n_11786, n_11787, n_11788, n_11789,
       n_11790;
  wire n_11791, n_11792, n_11793, n_11794, n_11795, n_11796, n_11797,
       n_11798;
  wire n_11799, n_11800, n_11801, n_11802, n_11803, n_11804, n_11805,
       n_11806;
  wire n_11807, n_11808, n_11809, n_11810, n_11811, n_11812, n_11813,
       n_11814;
  wire n_11815, n_11816, n_11817, n_11818, n_11819, n_11820, n_11821,
       n_11822;
  wire n_11823, n_11824, n_11825, n_11826, n_11827, n_11828, n_11829,
       n_11830;
  wire n_11831, n_11833, n_11834, n_11836, n_11838, n_11840, n_11842,
       n_11843;
  wire n_11844, n_11845, n_11846, n_11847, n_11848, n_11849, n_11850,
       n_11851;
  wire n_11852, n_11853, n_11854, n_11855, n_11856, n_11857, n_11858,
       n_11859;
  wire n_11860, n_11861, n_11862, n_11863, n_13034, n_14409_BAR,
       n_59812_BAR, n_61756_BAR;
  wire n_61758_BAR, n_61760_BAR, n_61762_BAR, n_61784_BAR, n_61792_BAR,
       n_61798_BAR, n_61804_BAR, n_61806_BAR;
  wire pcpi_div_wait, pcpi_div_wr, pcpi_mul_wr, pcpi_timeout,
       prefetched_high_word, \reg_op1[1]_9638 , \reg_op1[2]_9639 ,
       \reg_op1[3]_9640 ;
  wire \reg_op1[4]_9641 , \reg_op1[5]_9642 , \reg_op1[6]_9643 ,
       \reg_op1[7]_9644 , \reg_op1[8]_9645 , \reg_op1[9]_9646 ,
       \reg_op1[10]_9647 , \reg_op1[11]_9648 ;
  wire \reg_op1[12]_9649 , \reg_op1[13]_9650 , \reg_op1[14]_9651 ,
       \reg_op1[15]_9652 , \reg_op1[16]_9653 , \reg_op1[17]_9654 ,
       \reg_op1[18]_9655 , \reg_op1[19]_9656 ;
  wire \reg_op1[20]_9657 , \reg_op1[21]_9658 , \reg_op1[22]_9659 ,
       \reg_op1[23]_9660 , \reg_op1[24]_9661 , \reg_op1[25]_9662 ,
       \reg_op1[26]_9663 , \reg_op1[27]_9664 ;
  wire \reg_op1[28]_9665 , \reg_op1[29]_9666 , \reg_op1[30]_9667 ,
       \reg_op1[31]_9668 , \reg_op2[0]_9669 , \reg_op2[1]_9670 ,
       \reg_op2[2]_9671 , \reg_op2[3]_9672 ;
  wire \reg_op2[4]_9673 , \reg_op2[5]_9674 , \reg_op2[6]_9675 ,
       \reg_op2[7]_9676 , \reg_op2[8]_9677 , \reg_op2[9]_9678 ,
       \reg_op2[10]_9679 , \reg_op2[11]_9680 ;
  wire \reg_op2[12]_9681 , \reg_op2[13]_9682 , \reg_op2[14]_9683 ,
       \reg_op2[15]_9684 , \reg_op2[16]_9685 , \reg_op2[17]_9686 ,
       \reg_op2[18]_9687 , \reg_op2[19]_9688 ;
  wire \reg_op2[20]_9689 , \reg_op2[21]_9690 , \reg_op2[22]_9691 ,
       \reg_op2[23]_9692 , \reg_op2[24]_9693 , \reg_op2[25]_9694 ,
       \reg_op2[26]_9695 , \reg_op2[27]_9696 ;
  wire \reg_op2[28]_9697 , \reg_op2[29]_9698 , \reg_op2[30]_9699 ,
       \reg_op2[31]_9700 , sub_1235_38_Y_add_1235_58_n_1346,
       sub_1235_38_Y_add_1235_58_n_1348,
       sub_1235_38_Y_add_1235_58_n_1350,
       sub_1235_38_Y_add_1235_58_n_1352;
  wire sub_1235_38_Y_add_1235_58_n_1354,
       sub_1235_38_Y_add_1235_58_n_1356,
       sub_1235_38_Y_add_1235_58_n_1358,
       sub_1235_38_Y_add_1235_58_n_1360,
       sub_1235_38_Y_add_1235_58_n_1362,
       sub_1235_38_Y_add_1235_58_n_1364,
       sub_1235_38_Y_add_1235_58_n_1366,
       sub_1235_38_Y_add_1235_58_n_1368;
  wire sub_1235_38_Y_add_1235_58_n_1370,
       sub_1235_38_Y_add_1235_58_n_1372,
       sub_1235_38_Y_add_1235_58_n_1374,
       sub_1235_38_Y_add_1235_58_n_1376,
       sub_1235_38_Y_add_1235_58_n_1378,
       sub_1235_38_Y_add_1235_58_n_1380,
       sub_1235_38_Y_add_1235_58_n_1382,
       sub_1235_38_Y_add_1235_58_n_1384;
  wire sub_1235_38_Y_add_1235_58_n_1386,
       sub_1235_38_Y_add_1235_58_n_1388,
       sub_1235_38_Y_add_1235_58_n_1390,
       sub_1235_38_Y_add_1235_58_n_1392,
       sub_1235_38_Y_add_1235_58_n_1394,
       sub_1235_38_Y_add_1235_58_n_1396,
       sub_1235_38_Y_add_1235_58_n_1398,
       sub_1235_38_Y_add_1235_58_n_1400;
  wire sub_1235_38_Y_add_1235_58_n_1402,
       sub_1235_38_Y_add_1235_58_n_1404,
       sub_1235_38_Y_add_1235_58_n_1406,
       sub_1235_38_Y_add_1235_58_n_1407,
       sub_1235_38_Y_add_1235_58_n_1408,
       sub_1235_38_Y_add_1235_58_n_1410,
       sub_1235_38_Y_add_1235_58_n_1412,
       sub_1235_38_Y_add_1235_58_n_1413;
  wire sub_1235_38_Y_add_1235_58_n_1414,
       sub_1235_38_Y_add_1235_58_n_1415,
       sub_1235_38_Y_add_1235_58_n_1416,
       sub_1235_38_Y_add_1235_58_n_1417,
       sub_1235_38_Y_add_1235_58_n_1418,
       sub_1235_38_Y_add_1235_58_n_1419,
       sub_1235_38_Y_add_1235_58_n_1420,
       sub_1235_38_Y_add_1235_58_n_1421;
  wire sub_1235_38_Y_add_1235_58_n_1422,
       sub_1235_38_Y_add_1235_58_n_1423,
       sub_1235_38_Y_add_1235_58_n_1424,
       sub_1235_38_Y_add_1235_58_n_1425,
       sub_1235_38_Y_add_1235_58_n_1426,
       sub_1235_38_Y_add_1235_58_n_1427,
       sub_1235_38_Y_add_1235_58_n_1428,
       sub_1235_38_Y_add_1235_58_n_1429;
  wire sub_1235_38_Y_add_1235_58_n_1430,
       sub_1235_38_Y_add_1235_58_n_1431,
       sub_1235_38_Y_add_1235_58_n_1432,
       sub_1235_38_Y_add_1235_58_n_1433,
       sub_1235_38_Y_add_1235_58_n_1434,
       sub_1235_38_Y_add_1235_58_n_1435,
       sub_1235_38_Y_add_1235_58_n_1436,
       sub_1235_38_Y_add_1235_58_n_1437;
  wire sub_1235_38_Y_add_1235_58_n_1438,
       sub_1235_38_Y_add_1235_58_n_1439,
       sub_1235_38_Y_add_1235_58_n_1440,
       sub_1235_38_Y_add_1235_58_n_1441,
       sub_1235_38_Y_add_1235_58_n_1443;
  assign trace_data[0] = 1'b0;
  assign trace_data[1] = 1'b0;
  assign trace_data[2] = 1'b0;
  assign trace_data[3] = 1'b0;
  assign trace_data[4] = 1'b0;
  assign trace_data[5] = 1'b0;
  assign trace_data[6] = 1'b0;
  assign trace_data[7] = 1'b0;
  assign trace_data[8] = 1'b0;
  assign trace_data[9] = 1'b0;
  assign trace_data[10] = 1'b0;
  assign trace_data[11] = 1'b0;
  assign trace_data[12] = 1'b0;
  assign trace_data[13] = 1'b0;
  assign trace_data[14] = 1'b0;
  assign trace_data[15] = 1'b0;
  assign trace_data[16] = 1'b0;
  assign trace_data[17] = 1'b0;
  assign trace_data[18] = 1'b0;
  assign trace_data[19] = 1'b0;
  assign trace_data[20] = 1'b0;
  assign trace_data[21] = 1'b0;
  assign trace_data[22] = 1'b0;
  assign trace_data[23] = 1'b0;
  assign trace_data[24] = 1'b0;
  assign trace_data[25] = 1'b0;
  assign trace_data[26] = 1'b0;
  assign trace_data[27] = 1'b0;
  assign trace_data[28] = 1'b0;
  assign trace_data[29] = 1'b0;
  assign trace_data[30] = 1'b0;
  assign trace_data[31] = 1'b0;
  assign trace_data[32] = 1'b0;
  assign trace_data[33] = 1'b0;
  assign trace_data[34] = 1'b0;
  assign trace_data[35] = 1'b0;
  assign trace_valid = 1'b0;
  assign eoi[0] = 1'b0;
  assign eoi[1] = 1'b0;
  assign eoi[2] = 1'b0;
  assign eoi[3] = 1'b0;
  assign eoi[4] = 1'b0;
  assign eoi[5] = 1'b0;
  assign eoi[6] = 1'b0;
  assign eoi[7] = 1'b0;
  assign eoi[8] = 1'b0;
  assign eoi[9] = 1'b0;
  assign eoi[10] = 1'b0;
  assign eoi[11] = 1'b0;
  assign eoi[12] = 1'b0;
  assign eoi[13] = 1'b0;
  assign eoi[14] = 1'b0;
  assign eoi[15] = 1'b0;
  assign eoi[16] = 1'b0;
  assign eoi[17] = 1'b0;
  assign eoi[18] = 1'b0;
  assign eoi[19] = 1'b0;
  assign eoi[20] = 1'b0;
  assign eoi[21] = 1'b0;
  assign eoi[22] = 1'b0;
  assign eoi[23] = 1'b0;
  assign eoi[24] = 1'b0;
  assign eoi[25] = 1'b0;
  assign eoi[26] = 1'b0;
  assign eoi[27] = 1'b0;
  assign eoi[28] = 1'b0;
  assign eoi[29] = 1'b0;
  assign eoi[30] = 1'b0;
  assign eoi[31] = 1'b0;
  assign mem_la_addr[0] = 1'b0;
  assign mem_la_addr[1] = 1'b0;
  assign mem_addr[0] = 1'b0;
  assign mem_addr[1] = 1'b0;
  INVX20 g81907(.A (n_60), .Y (mem_la_write));
  INVX20 g81905(.A (n_150), .Y (mem_la_read));
  MX2X1 g82691__8428(.A (\genblk2.pcpi_div_dividend [0]), .B
       (\genblk2.pcpi_div_quotient [0]), .S0 (\genblk2.pcpi_div_n_2109
       ), .Y (\genblk2.pcpi_div_n_578 ));
  MX2X1 g82692__5526(.A (\genblk2.pcpi_div_dividend [30]), .B
       (\genblk2.pcpi_div_quotient [30]), .S0 (\genblk2.pcpi_div_n_2109
       ), .Y (\genblk2.pcpi_div_n_2111 ));
  MX2X1 g82694__3680(.A (\genblk2.pcpi_div_dividend [25]), .B
       (\genblk2.pcpi_div_quotient [25]), .S0 (\genblk2.pcpi_div_n_2109
       ), .Y (\genblk2.pcpi_div_n_2116 ));
  MX2X1 g82695__1617(.A (\genblk2.pcpi_div_dividend [19]), .B
       (\genblk2.pcpi_div_quotient [19]), .S0 (\genblk2.pcpi_div_n_2109
       ), .Y (\genblk2.pcpi_div_n_2122 ));
  MX2X1 g82697__1705(.A (\genblk2.pcpi_div_dividend [5]), .B
       (\genblk2.pcpi_div_quotient [5]), .S0 (\genblk2.pcpi_div_n_2109
       ), .Y (\genblk2.pcpi_div_n_2136 ));
  MX2X1 g82701__6131(.A (\genblk2.pcpi_div_dividend [17]), .B
       (\genblk2.pcpi_div_quotient [17]), .S0 (\genblk2.pcpi_div_n_2109
       ), .Y (\genblk2.pcpi_div_n_2124 ));
  MX2X1 g82702__1881(.A (\genblk2.pcpi_div_dividend [3]), .B
       (\genblk2.pcpi_div_quotient [3]), .S0 (\genblk2.pcpi_div_n_2109
       ), .Y (\genblk2.pcpi_div_n_2138 ));
  MX2X1 g82705__4733(.A (\genblk2.pcpi_div_dividend [1]), .B
       (\genblk2.pcpi_div_quotient [1]), .S0 (\genblk2.pcpi_div_n_2109
       ), .Y (\genblk2.pcpi_div_n_2140 ));
  MX2X1 g82706__6161(.A (\genblk2.pcpi_div_dividend [31]), .B
       (\genblk2.pcpi_div_quotient [31]), .S0 (\genblk2.pcpi_div_n_2109
       ), .Y (\genblk2.pcpi_div_n_2110 ));
  MX2X1 g82707__9315(.A (\genblk2.pcpi_div_dividend [7]), .B
       (\genblk2.pcpi_div_quotient [7]), .S0 (\genblk2.pcpi_div_n_2109
       ), .Y (\genblk2.pcpi_div_n_2134 ));
  MX2X1 g82708__9945(.A (\genblk2.pcpi_div_dividend [15]), .B
       (\genblk2.pcpi_div_quotient [15]), .S0 (\genblk2.pcpi_div_n_2109
       ), .Y (\genblk2.pcpi_div_n_2126 ));
  MX2X1 g82710__2346(.A (\genblk2.pcpi_div_dividend [13]), .B
       (\genblk2.pcpi_div_quotient [13]), .S0 (\genblk2.pcpi_div_n_2109
       ), .Y (\genblk2.pcpi_div_n_2128 ));
  MX2X1 g82711__1666(.A (\genblk2.pcpi_div_dividend [29]), .B
       (\genblk2.pcpi_div_quotient [29]), .S0 (\genblk2.pcpi_div_n_2109
       ), .Y (\genblk2.pcpi_div_n_2112 ));
  MX2X1 g82712__7410(.A (\genblk2.pcpi_div_dividend [27]), .B
       (\genblk2.pcpi_div_quotient [27]), .S0 (\genblk2.pcpi_div_n_2109
       ), .Y (\genblk2.pcpi_div_n_2114 ));
  MX2X1 g82715__2398(.A (\genblk2.pcpi_div_dividend [21]), .B
       (\genblk2.pcpi_div_quotient [21]), .S0 (\genblk2.pcpi_div_n_2109
       ), .Y (\genblk2.pcpi_div_n_2120 ));
  MX2X1 g82716__5107(.A (\genblk2.pcpi_div_dividend [11]), .B
       (\genblk2.pcpi_div_quotient [11]), .S0 (\genblk2.pcpi_div_n_2109
       ), .Y (\genblk2.pcpi_div_n_2130 ));
  MX2X1 g82720__5526(.A (\genblk2.pcpi_div_dividend [9]), .B
       (\genblk2.pcpi_div_quotient [9]), .S0 (\genblk2.pcpi_div_n_2109
       ), .Y (\genblk2.pcpi_div_n_2132 ));
  MX2X1 g82722__3680(.A (\genblk2.pcpi_div_dividend [23]), .B
       (\genblk2.pcpi_div_quotient [23]), .S0 (\genblk2.pcpi_div_n_2109
       ), .Y (\genblk2.pcpi_div_n_2118 ));
  OR2X2 g82723__1617(.A (\genblk2.pcpi_div_instr_div ), .B
       (\genblk2.pcpi_div_instr_divu ), .Y (\genblk2.pcpi_div_n_2109 ));
  DFFHQX1 \genblk2.pcpi_div_instr_divu_reg (.CK (clk), .D (n_6371), .Q
       (\genblk2.pcpi_div_instr_divu ));
  DFFHQX1 \genblk2.pcpi_div_instr_div_reg (.CK (clk), .D (n_6372), .Q
       (\genblk2.pcpi_div_instr_div ));
  NOR2BX1 g82726__2802(.AN (n_8138), .B (n_5597), .Y (n_6372));
  AND2X1 g82727__1705(.A (n_8138), .B (n_5597), .Y (n_6371));
  NAND4XL g82729__8246(.A (n_6369), .B (n_8325), .C (n_10451), .D
       (n_10551), .Y (n_6530));
  NOR4BX1 g82730__7098(.AN (resetn), .B (pcpi_div_wr), .C (n_5616), .D
       (n_6365), .Y (n_6369));
  NAND2XL g82734__7482(.A (n_5585), .B (n_5617), .Y (n_6365));
  DFFHQX1 \alu_out_q_reg[2] (.CK (clk), .D (n_6353), .Q (alu_out_q[2]));
  DFFHQX1 \alu_out_q_reg[3] (.CK (clk), .D (n_6352), .Q (alu_out_q[3]));
  DFFHQX1 \alu_out_q_reg[4] (.CK (clk), .D (n_6351), .Q (alu_out_q[4]));
  DFFHQX1 \alu_out_q_reg[5] (.CK (clk), .D (n_6350), .Q (alu_out_q[5]));
  DFFHQX1 \alu_out_q_reg[16] (.CK (clk), .D (n_6338), .Q
       (alu_out_q[16]));
  DFFHQX1 \alu_out_q_reg[17] (.CK (clk), .D (n_6349), .Q
       (alu_out_q[17]));
  DFFQXL \alu_out_q_reg[19] (.CK (clk), .D (n_6348), .Q
       (alu_out_q[19]));
  DFFQXL \alu_out_q_reg[20] (.CK (clk), .D (n_6347), .Q
       (alu_out_q[20]));
  DFFQXL \alu_out_q_reg[21] (.CK (clk), .D (n_6346), .Q
       (alu_out_q[21]));
  DFFQXL \alu_out_q_reg[22] (.CK (clk), .D (n_6345), .Q
       (alu_out_q[22]));
  DFFQXL \alu_out_q_reg[23] (.CK (clk), .D (n_6344), .Q
       (alu_out_q[23]));
  DFFQXL \alu_out_q_reg[24] (.CK (clk), .D (n_6337), .Q
       (alu_out_q[24]));
  DFFQXL \alu_out_q_reg[25] (.CK (clk), .D (n_6343), .Q
       (alu_out_q[25]));
  DFFQXL \alu_out_q_reg[26] (.CK (clk), .D (n_6342), .Q
       (alu_out_q[26]));
  DFFQXL \alu_out_q_reg[27] (.CK (clk), .D (n_6341), .Q
       (alu_out_q[27]));
  DFFQXL \alu_out_q_reg[28] (.CK (clk), .D (n_6336), .Q
       (alu_out_q[28]));
  DFFQXL \alu_out_q_reg[29] (.CK (clk), .D (n_6335), .Q
       (alu_out_q[29]));
  DFFQXL \alu_out_q_reg[30] (.CK (clk), .D (n_6340), .Q
       (alu_out_q[30]));
  DFFQXL \alu_out_q_reg[31] (.CK (clk), .D (n_6334), .Q
       (alu_out_q[31]));
  DFFRX1 decoder_pseudo_trigger_reg(.RN (1'b1), .CK (clk), .D (n_6307),
       .Q (UNCONNECTED), .QN (decoder_pseudo_trigger));
  DFFQXL \genblk1.pcpi_mul_rd_reg[0] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_91 ), .Q (\genblk1.pcpi_mul_rd [0]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[1] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_92 ), .Q (\genblk1.pcpi_mul_rd [1]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[2] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_93 ), .Q (\genblk1.pcpi_mul_rd [2]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[3] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_94 ), .Q (\genblk1.pcpi_mul_rd [3]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[4] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_95 ), .Q (\genblk1.pcpi_mul_rd [4]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[5] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_96 ), .Q (\genblk1.pcpi_mul_rd [5]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[6] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_97 ), .Q (\genblk1.pcpi_mul_rd [6]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[7] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_98 ), .Q (\genblk1.pcpi_mul_rd [7]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[8] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_99 ), .Q (\genblk1.pcpi_mul_rd [8]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[9] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_100 ), .Q (\genblk1.pcpi_mul_rd [9]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[10] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_101 ), .Q (\genblk1.pcpi_mul_rd [10]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[11] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_102 ), .Q (\genblk1.pcpi_mul_rd [11]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[12] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_103 ), .Q (\genblk1.pcpi_mul_rd [12]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[13] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_104 ), .Q (\genblk1.pcpi_mul_rd [13]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[14] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_105 ), .Q (\genblk1.pcpi_mul_rd [14]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[15] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_106 ), .Q (\genblk1.pcpi_mul_rd [15]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[16] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_107 ), .Q (\genblk1.pcpi_mul_rd [16]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[17] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_108 ), .Q (\genblk1.pcpi_mul_rd [17]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[18] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_109 ), .Q (\genblk1.pcpi_mul_rd [18]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[19] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_110 ), .Q (\genblk1.pcpi_mul_rd [19]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[20] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_111 ), .Q (\genblk1.pcpi_mul_rd [20]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[21] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_112 ), .Q (\genblk1.pcpi_mul_rd [21]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[22] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_113 ), .Q (\genblk1.pcpi_mul_rd [22]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[23] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_114 ), .Q (\genblk1.pcpi_mul_rd [23]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[24] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_115 ), .Q (\genblk1.pcpi_mul_rd [24]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[25] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_116 ), .Q (\genblk1.pcpi_mul_rd [25]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[26] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_117 ), .Q (\genblk1.pcpi_mul_rd [26]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[27] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_118 ), .Q (\genblk1.pcpi_mul_rd [27]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[28] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_119 ), .Q (\genblk1.pcpi_mul_rd [28]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[29] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_120 ), .Q (\genblk1.pcpi_mul_rd [29]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[30] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_121 ), .Q (\genblk1.pcpi_mul_rd [30]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[31] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_122 ), .Q (\genblk1.pcpi_mul_rd [31]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[32] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_123 ), .Q (\genblk1.pcpi_mul_rd [32]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[33] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_124 ), .Q (\genblk1.pcpi_mul_rd [33]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[34] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_125 ), .Q (\genblk1.pcpi_mul_rd [34]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[35] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_126 ), .Q (\genblk1.pcpi_mul_rd [35]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[36] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_127 ), .Q (\genblk1.pcpi_mul_rd [36]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[37] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_128 ), .Q (\genblk1.pcpi_mul_rd [37]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[38] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_129 ), .Q (\genblk1.pcpi_mul_rd [38]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[39] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_130 ), .Q (\genblk1.pcpi_mul_rd [39]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[40] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_131 ), .Q (\genblk1.pcpi_mul_rd [40]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[41] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_132 ), .Q (\genblk1.pcpi_mul_rd [41]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[42] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_133 ), .Q (\genblk1.pcpi_mul_rd [42]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[43] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_134 ), .Q (\genblk1.pcpi_mul_rd [43]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[44] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_135 ), .Q (\genblk1.pcpi_mul_rd [44]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[45] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_136 ), .Q (\genblk1.pcpi_mul_rd [45]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[46] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_137 ), .Q (\genblk1.pcpi_mul_rd [46]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[47] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_138 ), .Q (\genblk1.pcpi_mul_rd [47]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[48] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_139 ), .Q (\genblk1.pcpi_mul_rd [48]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[49] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_140 ), .Q (\genblk1.pcpi_mul_rd [49]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[50] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_141 ), .Q (\genblk1.pcpi_mul_rd [50]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[51] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_142 ), .Q (\genblk1.pcpi_mul_rd [51]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[52] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_143 ), .Q (\genblk1.pcpi_mul_rd [52]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[53] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_144 ), .Q (\genblk1.pcpi_mul_rd [53]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[54] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_145 ), .Q (\genblk1.pcpi_mul_rd [54]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[55] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_146 ), .Q (\genblk1.pcpi_mul_rd [55]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[56] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_147 ), .Q (\genblk1.pcpi_mul_rd [56]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[57] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_148 ), .Q (\genblk1.pcpi_mul_rd [57]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[58] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_149 ), .Q (\genblk1.pcpi_mul_rd [58]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[59] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_150 ), .Q (\genblk1.pcpi_mul_rd [59]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[60] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_151 ), .Q (\genblk1.pcpi_mul_rd [60]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[61] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_152 ), .Q (\genblk1.pcpi_mul_rd [61]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[62] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_153 ), .Q (\genblk1.pcpi_mul_rd [62]));
  DFFQXL \genblk1.pcpi_mul_rd_reg[63] (.CK (clk), .D
       (\genblk1.pcpi_mul_n_154 ), .Q (\genblk1.pcpi_mul_rd [63]));
  DFFQXL \genblk1.pcpi_mul_shift_out_reg (.CK (clk), .D (n_6285), .Q
       (\genblk1.pcpi_mul_shift_out ));
  DFFQXL \genblk2.pcpi_div_instr_rem_reg (.CK (clk), .D (n_6224), .Q
       (\genblk2.pcpi_div_instr_rem ));
  DFFQXL \genblk2.pcpi_div_instr_remu_reg (.CK (clk), .D (n_6223), .Q
       (\genblk2.pcpi_div_instr_remu ));
  DFFQXL \genblk2.pcpi_div_pcpi_rd_reg[0] (.CK (clk), .D
       (\genblk2.pcpi_div_n_578 ), .Q (pcpi_div_rd[0]));
  DFFQXL \genblk2.pcpi_div_pcpi_rd_reg[1] (.CK (clk), .D (n_6258), .Q
       (pcpi_div_rd[1]));
  DFFQXL \genblk2.pcpi_div_pcpi_rd_reg[2] (.CK (clk), .D (n_6257), .Q
       (pcpi_div_rd[2]));
  DFFQXL \genblk2.pcpi_div_pcpi_rd_reg[3] (.CK (clk), .D (n_6256), .Q
       (pcpi_div_rd[3]));
  DFFQXL \genblk2.pcpi_div_pcpi_rd_reg[4] (.CK (clk), .D (n_6255), .Q
       (pcpi_div_rd[4]));
  DFFQXL \genblk2.pcpi_div_pcpi_rd_reg[5] (.CK (clk), .D (n_6254), .Q
       (pcpi_div_rd[5]));
  DFFQXL \genblk2.pcpi_div_pcpi_rd_reg[6] (.CK (clk), .D (n_6253), .Q
       (pcpi_div_rd[6]));
  DFFQXL \genblk2.pcpi_div_pcpi_rd_reg[7] (.CK (clk), .D (n_6252), .Q
       (pcpi_div_rd[7]));
  DFFQXL \genblk2.pcpi_div_pcpi_rd_reg[8] (.CK (clk), .D (n_6251), .Q
       (pcpi_div_rd[8]));
  DFFQXL \genblk2.pcpi_div_pcpi_rd_reg[9] (.CK (clk), .D (n_6250), .Q
       (pcpi_div_rd[9]));
  DFFQXL \genblk2.pcpi_div_pcpi_rd_reg[10] (.CK (clk), .D (n_6249), .Q
       (pcpi_div_rd[10]));
  DFFQXL \genblk2.pcpi_div_pcpi_rd_reg[11] (.CK (clk), .D (n_6248), .Q
       (pcpi_div_rd[11]));
  DFFQXL \genblk2.pcpi_div_pcpi_rd_reg[12] (.CK (clk), .D (n_6247), .Q
       (pcpi_div_rd[12]));
  DFFQXL \genblk2.pcpi_div_pcpi_rd_reg[13] (.CK (clk), .D (n_6246), .Q
       (pcpi_div_rd[13]));
  DFFQXL \genblk2.pcpi_div_pcpi_rd_reg[14] (.CK (clk), .D (n_6245), .Q
       (pcpi_div_rd[14]));
  DFFQXL \genblk2.pcpi_div_pcpi_rd_reg[15] (.CK (clk), .D (n_6278), .Q
       (pcpi_div_rd[15]));
  DFFQXL \genblk2.pcpi_div_pcpi_rd_reg[16] (.CK (clk), .D (n_6244), .Q
       (pcpi_div_rd[16]));
  DFFQXL \genblk2.pcpi_div_pcpi_rd_reg[17] (.CK (clk), .D (n_6259), .Q
       (pcpi_div_rd[17]));
  DFFQXL \genblk2.pcpi_div_pcpi_rd_reg[18] (.CK (clk), .D (n_6243), .Q
       (pcpi_div_rd[18]));
  DFFQXL \genblk2.pcpi_div_pcpi_rd_reg[19] (.CK (clk), .D (n_6242), .Q
       (pcpi_div_rd[19]));
  DFFQXL \genblk2.pcpi_div_pcpi_rd_reg[20] (.CK (clk), .D (n_6241), .Q
       (pcpi_div_rd[20]));
  DFFQXL \genblk2.pcpi_div_pcpi_rd_reg[21] (.CK (clk), .D (n_6240), .Q
       (pcpi_div_rd[21]));
  DFFQXL \genblk2.pcpi_div_pcpi_rd_reg[22] (.CK (clk), .D (n_6239), .Q
       (pcpi_div_rd[22]));
  DFFQXL \genblk2.pcpi_div_pcpi_rd_reg[23] (.CK (clk), .D (n_6230), .Q
       (pcpi_div_rd[23]));
  DFFQXL \genblk2.pcpi_div_pcpi_rd_reg[24] (.CK (clk), .D (n_6238), .Q
       (pcpi_div_rd[24]));
  DFFQXL \genblk2.pcpi_div_pcpi_rd_reg[25] (.CK (clk), .D (n_6237), .Q
       (pcpi_div_rd[25]));
  DFFQXL \genblk2.pcpi_div_pcpi_rd_reg[26] (.CK (clk), .D (n_6236), .Q
       (pcpi_div_rd[26]));
  DFFQXL \genblk2.pcpi_div_pcpi_rd_reg[27] (.CK (clk), .D (n_6235), .Q
       (pcpi_div_rd[27]));
  DFFQXL \genblk2.pcpi_div_pcpi_rd_reg[28] (.CK (clk), .D (n_6234), .Q
       (pcpi_div_rd[28]));
  DFFQXL \genblk2.pcpi_div_pcpi_rd_reg[29] (.CK (clk), .D (n_6233), .Q
       (pcpi_div_rd[29]));
  DFFQXL \genblk2.pcpi_div_pcpi_rd_reg[30] (.CK (clk), .D (n_6232), .Q
       (pcpi_div_rd[30]));
  DFFQXL \genblk2.pcpi_div_pcpi_rd_reg[31] (.CK (clk), .D (n_6231), .Q
       (pcpi_div_rd[31]));
  DFFHQX1 \genblk2.pcpi_div_pcpi_wait_q_reg (.CK (clk), .D (n_6293), .Q
       (\genblk2.pcpi_div_pcpi_wait_q ));
  DFFQXL is_compare_reg(.CK (clk), .D (n_6311), .Q (is_compare));
  DFFQXL is_lbu_lhu_lw_reg(.CK (clk), .D (n_6095), .Q (is_lbu_lhu_lw));
  DFFQX2 is_lui_auipc_jal_jalr_addi_add_sub_reg(.CK (clk), .D (n_6312),
       .Q (is_lui_auipc_jal_jalr_addi_add_sub));
  DFFHQX1 is_lui_auipc_jal_reg(.CK (clk), .D (n_6085), .Q
       (is_lui_auipc_jal));
  DFFQXL is_slti_blt_slt_reg(.CK (clk), .D (n_6086), .Q
       (is_slti_blt_slt));
  DFFQXL is_sltiu_bltu_sltu_reg(.CK (clk), .D (n_6127), .Q
       (is_sltiu_bltu_sltu));
  DFFHQX1 last_mem_valid_reg(.CK (clk), .D (n_6068), .Q
       (last_mem_valid));
  DFFHQX1 pcpi_timeout_reg(.CK (clk), .D (n_6274), .Q (pcpi_timeout));
  DFFQXL \reg_out_reg[0] (.CK (clk), .D (n_6339), .Q (reg_out[0]));
  OAI2BB1X1 g89561__4733(.A0N (n_5997), .A1N (n_208), .B0 (n_6133), .Y
       (current_pc[27]));
  OAI2BB1X1 g89562__6161(.A0N (n_5997), .A1N (n_214), .B0 (n_6138), .Y
       (current_pc[30]));
  OAI2BB1X1 g89563__9315(.A0N (n_5997), .A1N (n_164), .B0 (n_6149), .Y
       (current_pc[5]));
  OAI2BB1X1 g89564__9945(.A0N (n_5997), .A1N (n_170), .B0 (n_6150), .Y
       (current_pc[4]));
  OAI2BB1X1 g89565__2883(.A0N (n_168), .A1N (n_5997), .B0 (n_6151), .Y
       (current_pc[3]));
  OAI2BB1X1 g89566__2346(.A0N (n_166), .A1N (n_5997), .B0 (n_6152), .Y
       (current_pc[2]));
  OAI2BB1X1 g89567__1666(.A0N (n_5997), .A1N (n_212), .B0 (n_6135), .Y
       (current_pc[29]));
  OAI2BB1X1 g89568__7410(.A0N (n_5997), .A1N (n_210), .B0 (n_6148), .Y
       (current_pc[28]));
  OAI2BB1X1 g89569__6417(.A0N (n_5997), .A1N (n_216), .B0 (n_6145), .Y
       (current_pc[31]));
  OAI2BB1X1 g89570__5477(.A0N (n_5997), .A1N (n_206), .B0 (n_6131), .Y
       (current_pc[26]));
  OAI2BB1X1 g89571__2398(.A0N (n_5997), .A1N (n_204), .B0 (n_6129), .Y
       (current_pc[25]));
  OAI2BB1X1 g89572__5107(.A0N (n_5997), .A1N (n_202), .B0 (n_6128), .Y
       (current_pc[24]));
  OAI2BB1X1 g89573__6260(.A0N (n_5997), .A1N (n_200), .B0 (n_6100), .Y
       (current_pc[23]));
  OAI2BB1X1 g89574__4319(.A0N (n_5997), .A1N (n_146), .B0 (n_6093), .Y
       (current_pc[22]));
  OAI2BB1X1 g89575__8428(.A0N (n_5997), .A1N (n_144), .B0 (n_6102), .Y
       (current_pc[21]));
  OAI2BB1X1 g89576__5526(.A0N (n_5997), .A1N (n_198), .B0 (n_6099), .Y
       (current_pc[20]));
  OAI2BB1X1 g89577__6783(.A0N (n_5997), .A1N (n_142), .B0 (n_6089), .Y
       (current_pc[19]));
  OAI2BB1X1 g89578__3680(.A0N (n_5997), .A1N (n_194), .B0 (n_6084), .Y
       (current_pc[17]));
  OAI2BB1X1 g89579__1617(.A0N (n_5997), .A1N (n_192), .B0 (n_6083), .Y
       (current_pc[16]));
  MX2X1 g89580__2802(.A (reg_out[27]), .B (alu_out_q[27]), .S0
       (latched_stalu), .Y (n_208));
  MX2X1 g89581__1705(.A (reg_out[4]), .B (alu_out_q[4]), .S0
       (latched_stalu), .Y (n_170));
  MX2X1 g89582__5122(.A (reg_out[3]), .B (alu_out_q[3]), .S0
       (latched_stalu), .Y (n_168));
  MX2X1 g89583__8246(.A (reg_out[2]), .B (alu_out_q[2]), .S0
       (latched_stalu), .Y (n_166));
  MX2X1 g89584__7098(.A (reg_out[31]), .B (alu_out_q[31]), .S0
       (latched_stalu), .Y (n_216));
  MX2X1 g89585__6131(.A (reg_out[30]), .B (alu_out_q[30]), .S0
       (latched_stalu), .Y (n_214));
  MX2X1 g89586__1881(.A (reg_out[29]), .B (alu_out_q[29]), .S0
       (latched_stalu), .Y (n_212));
  MX2X1 g89587__5115(.A (reg_out[28]), .B (alu_out_q[28]), .S0
       (latched_stalu), .Y (n_210));
  MX2X1 g89588__7482(.A (reg_out[5]), .B (alu_out_q[5]), .S0
       (latched_stalu), .Y (n_164));
  MX2X1 g89589__4733(.A (reg_out[25]), .B (alu_out_q[25]), .S0
       (latched_stalu), .Y (n_204));
  MX2X1 g89590__6161(.A (reg_out[26]), .B (alu_out_q[26]), .S0
       (latched_stalu), .Y (n_206));
  MX2X1 g89591__9315(.A (reg_out[24]), .B (alu_out_q[24]), .S0
       (latched_stalu), .Y (n_202));
  MX2X1 g89592__9945(.A (reg_out[23]), .B (alu_out_q[23]), .S0
       (latched_stalu), .Y (n_200));
  MX2X1 g89593__2883(.A (reg_out[22]), .B (alu_out_q[22]), .S0
       (latched_stalu), .Y (n_146));
  MX2X1 g89594__2346(.A (reg_out[21]), .B (alu_out_q[21]), .S0
       (latched_stalu), .Y (n_144));
  MX2X1 g89595__1666(.A (reg_out[20]), .B (alu_out_q[20]), .S0
       (latched_stalu), .Y (n_198));
  MX2X1 g89596__7410(.A (reg_out[19]), .B (alu_out_q[19]), .S0
       (latched_stalu), .Y (n_142));
  MX2X1 g89597__6417(.A (reg_out[17]), .B (alu_out_q[17]), .S0
       (latched_stalu), .Y (n_194));
  MX2X1 g89598__5477(.A (reg_out[16]), .B (alu_out_q[16]), .S0
       (latched_stalu), .Y (n_192));
  OAI211X1 g89619__2398(.A0 (n_6035), .A1 (n_119), .B0 (n_6220), .C0
       (n_6331), .Y (n_6353));
  OAI211X1 g89620__5107(.A0 (n_6037), .A1 (n_119), .B0 (n_6219), .C0
       (n_6330), .Y (n_6352));
  OAI211X1 g89621__6260(.A0 (n_6028), .A1 (n_119), .B0 (n_6218), .C0
       (n_6329), .Y (n_6351));
  OAI211X1 g89622__4319(.A0 (n_6055), .A1 (n_119), .B0 (n_6217), .C0
       (n_6328), .Y (n_6350));
  OAI221X1 g89623__8428(.A0 (n_278), .A1 (n_6088), .B0 (n_6056), .B1
       (n_119), .C0 (n_6326), .Y (n_6349));
  OAI211X1 g89624__5526(.A0 (n_6040), .A1 (n_119), .B0 (n_6216), .C0
       (n_6325), .Y (n_6348));
  OAI221X1 g89625__6783(.A0 (n_278), .A1 (n_6090), .B0 (n_6030), .B1
       (n_119), .C0 (n_6324), .Y (n_6347));
  OAI211X1 g89626__3680(.A0 (n_6039), .A1 (n_119), .B0 (n_6215), .C0
       (n_6321), .Y (n_6346));
  OAI211X1 g89627__1617(.A0 (n_6054), .A1 (n_119), .B0 (n_6214), .C0
       (n_6323), .Y (n_6345));
  OAI211X1 g89628__2802(.A0 (n_6031), .A1 (n_119), .B0 (n_6213), .C0
       (n_6322), .Y (n_6344));
  OAI221X1 g89629__1705(.A0 (n_278), .A1 (n_6091), .B0 (n_6038), .B1
       (n_119), .C0 (n_6319), .Y (n_6343));
  OAI221X1 g89630__5122(.A0 (n_278), .A1 (n_6092), .B0 (n_6033), .B1
       (n_119), .C0 (n_6318), .Y (n_6342));
  OAI211X1 g89631__8246(.A0 (n_6041), .A1 (n_119), .B0 (n_6212), .C0
       (n_6317), .Y (n_6341));
  OAI211X1 g89632__7098(.A0 (n_6036), .A1 (n_119), .B0 (n_6211), .C0
       (n_6314), .Y (n_6340));
  NAND2X1 g89633__6131(.A (n_6294), .B (n_6332), .Y (n_6339));
  OAI211X1 g89634__1881(.A0 (n_6053), .A1 (n_119), .B0 (n_6273), .C0
       (n_6327), .Y (n_6338));
  OAI211X1 g89635__5115(.A0 (n_6032), .A1 (n_119), .B0 (n_6272), .C0
       (n_6320), .Y (n_6337));
  OAI211X1 g89636__7482(.A0 (n_6043), .A1 (n_119), .B0 (n_6271), .C0
       (n_6316), .Y (n_6336));
  OAI211X1 g89637__4733(.A0 (n_6044), .A1 (n_119), .B0 (n_6270), .C0
       (n_6315), .Y (n_6335));
  OAI221X1 g89638__6161(.A0 (n_6051), .A1 (n_119), .B0 (n_6059), .B1
       (n_6048), .C0 (n_6333), .Y (n_6334));
  AOI22XL g89639__9315(.A0 (is_lui_auipc_jal_jalr_addi_add_sub), .A1
       (n_6656), .B0 (n_279), .B1 (n_11691), .Y (n_6333));
  AOI22XL g89640__9945(.A0 (cpu_state[5]), .A1 (n_6313), .B0
       (decoded_imm[0]), .B1 (cpu_state[3]), .Y (n_6332));
  AOI32X1 g89641__2883(.A0 (\reg_op1[2]_9639 ), .A1 (\reg_op2[2]_9671
       ), .A2 (n_283), .B0 (is_lui_auipc_jal_jalr_addi_add_sub), .B1
       (n_6627), .Y (n_6331));
  AOI32X1 g89642__2346(.A0 (\reg_op1[3]_9640 ), .A1 (\reg_op2[3]_9672
       ), .A2 (n_283), .B0 (is_lui_auipc_jal_jalr_addi_add_sub), .B1
       (n_6628), .Y (n_6330));
  AOI32X1 g89643__1666(.A0 (\reg_op1[4]_9641 ), .A1 (\reg_op2[4]_9673
       ), .A2 (n_283), .B0 (is_lui_auipc_jal_jalr_addi_add_sub), .B1
       (n_6629), .Y (n_6329));
  AOI32X1 g89644__7410(.A0 (\reg_op1[5]_9642 ), .A1 (\reg_op2[5]_9674
       ), .A2 (n_283), .B0 (is_lui_auipc_jal_jalr_addi_add_sub), .B1
       (n_6630), .Y (n_6328));
  AOI32X1 g89645__6417(.A0 (\reg_op2[16]_9685 ), .A1 (\reg_op1[16]_9653
       ), .A2 (n_283), .B0 (is_lui_auipc_jal_jalr_addi_add_sub), .B1
       (n_6641), .Y (n_6327));
  AOI32X1 g89646__5477(.A0 (\reg_op2[17]_9686 ), .A1 (\reg_op1[17]_9654
       ), .A2 (n_283), .B0 (is_lui_auipc_jal_jalr_addi_add_sub), .B1
       (n_6642), .Y (n_6326));
  AOI32X1 g89647__2398(.A0 (\reg_op2[19]_9688 ), .A1 (\reg_op1[19]_9656
       ), .A2 (n_283), .B0 (is_lui_auipc_jal_jalr_addi_add_sub), .B1
       (n_6644), .Y (n_6325));
  AOI32X1 g89648__5107(.A0 (\reg_op2[20]_9689 ), .A1 (\reg_op1[20]_9657
       ), .A2 (n_283), .B0 (is_lui_auipc_jal_jalr_addi_add_sub), .B1
       (n_6645), .Y (n_6324));
  AOI32X1 g89649__6260(.A0 (\reg_op2[22]_9691 ), .A1 (\reg_op1[22]_9659
       ), .A2 (n_283), .B0 (is_lui_auipc_jal_jalr_addi_add_sub), .B1
       (n_6647), .Y (n_6323));
  AOI32X1 g89650__4319(.A0 (\reg_op2[23]_9692 ), .A1 (\reg_op1[23]_9660
       ), .A2 (n_283), .B0 (is_lui_auipc_jal_jalr_addi_add_sub), .B1
       (n_6648), .Y (n_6322));
  AOI32X1 g89651__8428(.A0 (\reg_op2[21]_9690 ), .A1 (\reg_op1[21]_9658
       ), .A2 (n_283), .B0 (is_lui_auipc_jal_jalr_addi_add_sub), .B1
       (n_6646), .Y (n_6321));
  AOI32X1 g89652__5526(.A0 (\reg_op2[24]_9693 ), .A1 (\reg_op1[24]_9661
       ), .A2 (n_283), .B0 (is_lui_auipc_jal_jalr_addi_add_sub), .B1
       (n_6649), .Y (n_6320));
  AOI32X1 g89653__6783(.A0 (\reg_op2[25]_9694 ), .A1 (\reg_op1[25]_9662
       ), .A2 (n_283), .B0 (is_lui_auipc_jal_jalr_addi_add_sub), .B1
       (n_6650), .Y (n_6319));
  AOI32X1 g89654__3680(.A0 (\reg_op2[26]_9695 ), .A1 (\reg_op1[26]_9663
       ), .A2 (n_283), .B0 (is_lui_auipc_jal_jalr_addi_add_sub), .B1
       (n_6651), .Y (n_6318));
  AOI32X1 g89655__1617(.A0 (\reg_op2[27]_9696 ), .A1 (\reg_op1[27]_9664
       ), .A2 (n_283), .B0 (is_lui_auipc_jal_jalr_addi_add_sub), .B1
       (n_6652), .Y (n_6317));
  AOI32X1 g89656__2802(.A0 (\reg_op2[28]_9697 ), .A1 (\reg_op1[28]_9665
       ), .A2 (n_283), .B0 (is_lui_auipc_jal_jalr_addi_add_sub), .B1
       (n_6653), .Y (n_6316));
  AOI32X1 g89657__1705(.A0 (\reg_op2[29]_9698 ), .A1 (\reg_op1[29]_9666
       ), .A2 (n_283), .B0 (is_lui_auipc_jal_jalr_addi_add_sub), .B1
       (n_6654), .Y (n_6315));
  AOI32X1 g89658__5122(.A0 (\reg_op2[30]_9699 ), .A1 (\reg_op1[30]_9667
       ), .A2 (n_283), .B0 (is_lui_auipc_jal_jalr_addi_add_sub), .B1
       (n_6655), .Y (n_6314));
  NAND4XL g89661__8246(.A (n_6067), .B (n_6066), .C (n_6309), .D
       (n_6310), .Y (n_6313));
  NOR2X1 g89662__7098(.A (n_538), .B (n_6227), .Y (n_6312));
  AOI21X1 g89663__6131(.A0 (n_6201), .A1 (n_130), .B0 (n_538), .Y
       (n_6311));
  AND2X4 g89664__1881(.A (decoder_pseudo_trigger), .B
       (decoder_trigger), .Y (n_538));
  AOI22XL g89665__5115(.A0 (\genblk1.pcpi_mul_rd [32]), .A1 (n_11690),
       .B0 (pcpi_rd[0]), .B1 (n_11689), .Y (n_6310));
  AOI22X1 g89666__7482(.A0 (\genblk1.pcpi_mul_rd [0]), .A1
       (n_59812_BAR), .B0 (pcpi_div_rd[0]), .B1 (n_39), .Y (n_6309));
  NOR2X4 g89668__4733(.A (\genblk1.pcpi_mul_shift_out ), .B (n_6527),
       .Y (n_59812_BAR));
  NOR3X1 g89670__6161(.A (mem_do_prefetch), .B (n_6063), .C (mem_done),
       .Y (n_6307));
  NAND2BXL g89673__9945(.AN (n_356), .B (pcpi_div_wr), .Y (n_40));
  NAND2BX1 g89676__2346(.AN (n_356), .B (pcpi_mul_wr), .Y (n_6527));
  NAND2X1 g89677__1666(.A (resetn), .B (n_6304), .Y (n_150));
  OAI211X1 g89678__7410(.A0 (n_6524), .A1 (n_6302), .B0 (resetn), .C0
       (n_6295), .Y (mem_done));
  NAND2X1 g89679__6417(.A (n_278), .B (n_6303), .Y (n_356));
  OAI32X1 g89680__5477(.A0 (mem_la_secondword), .A1 (n_6291), .A2
       (n_276), .B0 (n_158), .B1 (n_5970), .Y (n_6304));
  NOR4X1 g89681__2398(.A (instr_rdinstrh), .B (instr_rdinstr), .C
       (n_120), .D (n_6301), .Y (n_6303));
  NOR2BX1 g89682__5107(.AN (n_276), .B (n_6292), .Y (n_6302));
  MX2X1 g89691__1705(.A (reg_op1[0]), .B (\genblk2.pcpi_div_divisor
       [0]), .S0 (\genblk2.pcpi_div_n_4742 ), .Y
       (\genblk2.pcpi_div_n_1929 ));
  OR4X1 g89698__7482(.A (instr_rdcycleh), .B (instr_rdcycle), .C
       (n_6086), .D (n_6298), .Y (n_6301));
  NAND2X1 g89699__4733(.A (mem_rdata_latched[1]), .B
       (mem_rdata_latched[0]), .Y (n_276));
  AND2X1 g89718__2802(.A (\genblk2.pcpi_div_dividend [30]), .B
       (\genblk2.pcpi_div_n_4742 ), .Y (\genblk2.pcpi_div_n_1867 ));
  AND2X1 g89719__1705(.A (\genblk2.pcpi_div_dividend [29]), .B
       (\genblk2.pcpi_div_n_4742 ), .Y (\genblk2.pcpi_div_n_1868 ));
  AND2X1 g89720__5122(.A (\genblk2.pcpi_div_dividend [27]), .B
       (\genblk2.pcpi_div_n_4742 ), .Y (\genblk2.pcpi_div_n_1870 ));
  AND2X1 g89721__8246(.A (\genblk2.pcpi_div_dividend [28]), .B
       (\genblk2.pcpi_div_n_4742 ), .Y (\genblk2.pcpi_div_n_1869 ));
  AND2X1 g89722__7098(.A (\genblk2.pcpi_div_dividend [26]), .B
       (\genblk2.pcpi_div_n_4742 ), .Y (\genblk2.pcpi_div_n_1871 ));
  AND2X1 g89723__6131(.A (\genblk2.pcpi_div_dividend [25]), .B
       (\genblk2.pcpi_div_n_4742 ), .Y (\genblk2.pcpi_div_n_1872 ));
  AND2X1 g89724__1881(.A (\genblk2.pcpi_div_dividend [24]), .B
       (\genblk2.pcpi_div_n_4742 ), .Y (\genblk2.pcpi_div_n_1873 ));
  AND2X1 g89725__5115(.A (\genblk2.pcpi_div_dividend [23]), .B
       (\genblk2.pcpi_div_n_4742 ), .Y (\genblk2.pcpi_div_n_1874 ));
  AND2X1 g89726__7482(.A (\genblk2.pcpi_div_dividend [22]), .B
       (\genblk2.pcpi_div_n_4742 ), .Y (\genblk2.pcpi_div_n_1875 ));
  AND2X1 g89727__4733(.A (\genblk2.pcpi_div_dividend [21]), .B
       (\genblk2.pcpi_div_n_4742 ), .Y (\genblk2.pcpi_div_n_1876 ));
  AND2X1 g89728__6161(.A (\genblk2.pcpi_div_dividend [20]), .B
       (\genblk2.pcpi_div_n_4742 ), .Y (\genblk2.pcpi_div_n_1877 ));
  AND2X1 g89729__9315(.A (\genblk2.pcpi_div_dividend [19]), .B
       (\genblk2.pcpi_div_n_4742 ), .Y (\genblk2.pcpi_div_n_1878 ));
  AND2X1 g89730__9945(.A (\genblk2.pcpi_div_dividend [18]), .B
       (\genblk2.pcpi_div_n_4742 ), .Y (\genblk2.pcpi_div_n_1879 ));
  AND2X1 g89731__2883(.A (\genblk2.pcpi_div_dividend [17]), .B
       (\genblk2.pcpi_div_n_4742 ), .Y (\genblk2.pcpi_div_n_1880 ));
  AND2X1 g89732__2346(.A (\genblk2.pcpi_div_dividend [16]), .B
       (\genblk2.pcpi_div_n_4742 ), .Y (\genblk2.pcpi_div_n_1881 ));
  AND2X1 g89733__1666(.A (\genblk2.pcpi_div_dividend [15]), .B
       (\genblk2.pcpi_div_n_4742 ), .Y (\genblk2.pcpi_div_n_1882 ));
  AND2X1 g89734__7410(.A (\genblk2.pcpi_div_dividend [14]), .B
       (\genblk2.pcpi_div_n_4742 ), .Y (\genblk2.pcpi_div_n_1883 ));
  AND2X1 g89735__6417(.A (\genblk2.pcpi_div_dividend [13]), .B
       (\genblk2.pcpi_div_n_4742 ), .Y (\genblk2.pcpi_div_n_1884 ));
  AND2X1 g89736__5477(.A (\genblk2.pcpi_div_dividend [12]), .B
       (\genblk2.pcpi_div_n_4742 ), .Y (\genblk2.pcpi_div_n_1885 ));
  AND2X1 g89737__2398(.A (\genblk2.pcpi_div_dividend [11]), .B
       (\genblk2.pcpi_div_n_4742 ), .Y (\genblk2.pcpi_div_n_1886 ));
  AND2X1 g89738__5107(.A (\genblk2.pcpi_div_dividend [10]), .B
       (\genblk2.pcpi_div_n_4742 ), .Y (\genblk2.pcpi_div_n_1887 ));
  AND2X1 g89739__6260(.A (\genblk2.pcpi_div_dividend [9]), .B
       (\genblk2.pcpi_div_n_4742 ), .Y (\genblk2.pcpi_div_n_1888 ));
  AND2X1 g89740__4319(.A (\genblk2.pcpi_div_dividend [8]), .B
       (\genblk2.pcpi_div_n_4742 ), .Y (\genblk2.pcpi_div_n_1889 ));
  AND2X1 g89741__8428(.A (\genblk2.pcpi_div_dividend [7]), .B
       (\genblk2.pcpi_div_n_4742 ), .Y (\genblk2.pcpi_div_n_1890 ));
  AND2X1 g89742__5526(.A (\genblk2.pcpi_div_dividend [6]), .B
       (\genblk2.pcpi_div_n_4742 ), .Y (\genblk2.pcpi_div_n_1891 ));
  AND2X1 g89743__6783(.A (\genblk2.pcpi_div_dividend [5]), .B
       (\genblk2.pcpi_div_n_4742 ), .Y (\genblk2.pcpi_div_n_1892 ));
  AND2X1 g89744__3680(.A (\genblk2.pcpi_div_dividend [4]), .B
       (\genblk2.pcpi_div_n_4742 ), .Y (\genblk2.pcpi_div_n_1893 ));
  AND2X1 g89745__1617(.A (\genblk2.pcpi_div_dividend [3]), .B
       (\genblk2.pcpi_div_n_4742 ), .Y (\genblk2.pcpi_div_n_1894 ));
  AND2X1 g89746__2802(.A (\genblk2.pcpi_div_dividend [2]), .B
       (\genblk2.pcpi_div_n_4742 ), .Y (\genblk2.pcpi_div_n_1895 ));
  AND2X1 g89747__1705(.A (\genblk2.pcpi_div_dividend [1]), .B
       (\genblk2.pcpi_div_n_4742 ), .Y (\genblk2.pcpi_div_n_1896 ));
  AND2X1 g89748__5122(.A (\genblk2.pcpi_div_dividend [0]), .B
       (\genblk2.pcpi_div_n_4742 ), .Y (\genblk2.pcpi_div_n_1897 ));
  OAI211X1 g89749__8246(.A0 (n_6011), .A1 (n_46), .B0 (n_6296), .C0
       (n_6299), .Y (mem_rdata_latched[0]));
  OAI211X1 g89750__7098(.A0 (n_6027), .A1 (n_46), .B0 (n_6297), .C0
       (n_6300), .Y (mem_rdata_latched[1]));
  OR2X4 g89751__6131(.A (\genblk2.pcpi_div_pcpi_wait_q ), .B (n_5999),
       .Y (\genblk2.pcpi_div_n_4742 ));
  AOI22XL g89752__1881(.A0 (n_567), .A1 (n_6865), .B0
       (mem_16bit_buffer[1]), .B1 (n_360), .Y (n_6300));
  AOI22XL g89753__5115(.A0 (n_567), .A1 (n_6864), .B0
       (mem_16bit_buffer[0]), .B1 (n_360), .Y (n_6299));
  NAND4XL g89755__7482(.A (n_6042), .B (n_6061), .C (n_6227), .D
       (n_6288), .Y (n_6298));
  NAND2BXL g89756__4733(.AN (n_113), .B (mem_rdata_q[1]), .Y (n_6297));
  NAND2BXL g89757__6161(.AN (n_113), .B (mem_rdata_q[0]), .Y (n_6296));
  NAND2X1 g89758__9315(.A (n_6567), .B (n_6292), .Y (n_6295));
  AOI22XL g89759__9945(.A0 (cpu_state[0]), .A1 (n_6289), .B0
       (cpu_state[2]), .B1 (reg_op1[0]), .Y (n_6294));
  NOR2X1 g89760__2883(.A (n_5999), .B (n_544), .Y (n_6293));
  MX2X1 g89761__2346(.A (mem_rdata_q[17]), .B (mem_rdata[17]), .S0
       (mem_xfer), .Y (n_6865));
  MX2X1 g89762__1666(.A (mem_rdata_q[16]), .B (mem_rdata[16]), .S0
       (mem_xfer), .Y (n_6864));
  NAND2BX1 g89765__7410(.AN (n_268), .B (mem_xfer), .Y (n_46));
  INVX1 g89766(.A (mem_la_firstword_xfer), .Y (n_6291));
  OAI211X1 g89767__6417(.A0 (mem_do_rinst), .A1 (n_6555), .B0 (n_6050),
       .C0 (mem_xfer), .Y (n_6292));
  OAI22X1 g89768__5477(.A0 (n_6275), .A1 (n_6287), .B0 (n_6283), .B1
       (n_6060), .Y (mem_la_firstword_xfer));
  OR2X1 g89769__2398(.A (n_268), .B (mem_xfer), .Y (n_113));
  NOR2X1 g89772__5107(.A (n_6284), .B (n_544), .Y (n_6290));
  OAI211X1 g89773__6260(.A0 (n_343), .A1 (n_6011), .B0 (n_6276), .C0
       (n_6229), .Y (n_6289));
  NOR4X1 g89774__4319(.A (instr_sw), .B (instr_sh), .C (instr_bgeu), .D
       (n_6282), .Y (n_6288));
  INVX1 g89776(.A (n_567), .Y (n_277));
  NAND2X1 g89777__8428(.A (mem_do_rinst), .B (n_5970), .Y (n_6287));
  NOR2X1 g89778__5526(.A (n_6524), .B (n_5970), .Y (n_567));
  OR2X1 g89779__6783(.A (mem_la_secondword), .B (n_5970), .Y (n_360));
  AOI2BB1X1 g89780__3680(.A0N (n_5597), .A1N (n_5598), .B0 (n_6565), .Y
       (n_6285));
  NOR4X1 g89781__1617(.A (\genblk2.pcpi_div_instr_remu ), .B
       (\genblk2.pcpi_div_instr_rem ), .C (\genblk2.pcpi_div_instr_divu
       ), .D (\genblk2.pcpi_div_instr_div ), .Y (n_6284));
  MXI2XL g89782__2802(.A (n_6280), .B (mem_la_firstword_reg), .S0
       (last_mem_valid), .Y (n_6283));
  NAND3X1 g89783__1705(.A (n_6048), .B (n_6094), .C (n_6228), .Y
       (n_6282));
  OR2X1 g89784__5122(.A (mem_la_secondword), .B (n_6280), .Y (n_268));
  OR3X1 g89786__8246(.A (n_5599), .B (n_6260), .C (n_544), .Y (n_6565));
  INVX1 g89805(.A (n_6524), .Y (n_6280));
  NAND3BXL g89821__7098(.AN (n_340), .B (n_311), .C (n_331), .Y
       (n_343));
  NAND2X1 g89822__6131(.A (n_313), .B (n_6266), .Y (n_6524));
  OAI2BB1X1 g89824__5115(.A0N (\genblk2.pcpi_div_quotient [15]), .A1N
       (n_5694), .B0 (n_6179), .Y (n_6278));
  NAND2X1 g89826__4733(.A (n_340), .B (mem_rdata[16]), .Y (n_6276));
  NOR2BX1 g89827__6161(.AN (last_mem_valid), .B (mem_la_firstword_reg),
       .Y (n_6275));
  NOR2X1 g89828__9315(.A (n_258), .B (n_544), .Y (n_6274));
  NAND2X1 g89829__9945(.A (n_279), .B (n_6661), .Y (n_6273));
  NAND2X1 g89830__2883(.A (n_279), .B (n_6668), .Y (n_6272));
  NAND2X1 g89831__2346(.A (n_279), .B (n_6672), .Y (n_6271));
  NAND2X1 g89832__1666(.A (n_279), .B (n_6673), .Y (n_6270));
  NOR2X1 g89836__2398(.A (mem_la_secondword), .B (n_6160), .Y (n_6266));
  OAI2BB1X1 g89843__6783(.A0N (n_5997), .A1N (n_188), .B0 (n_6130), .Y
       (current_pc[14]));
  OAI2BB1X1 g89844__3680(.A0N (n_5997), .A1N (n_172), .B0 (n_6132), .Y
       (current_pc[13]));
  OAI2BB1X1 g89845__1617(.A0N (n_5997), .A1N (n_186), .B0 (n_6136), .Y
       (current_pc[12]));
  OAI2BB1X1 g89846__2802(.A0N (n_5997), .A1N (n_184), .B0 (n_6137), .Y
       (current_pc[11]));
  OAI2BB1X1 g89847__1705(.A0N (n_5997), .A1N (n_182), .B0 (n_6140), .Y
       (current_pc[10]));
  OAI2BB1X1 g89848__5122(.A0N (n_5997), .A1N (n_180), .B0 (n_6142), .Y
       (current_pc[9]));
  OAI2BB1X1 g89849__8246(.A0N (n_5997), .A1N (n_178), .B0 (n_6143), .Y
       (current_pc[8]));
  OAI2BB1X1 g89850__7098(.A0N (n_5997), .A1N (n_176), .B0 (n_6144), .Y
       (current_pc[7]));
  OAI2BB1X1 g89851__6131(.A0N (n_5997), .A1N (n_174), .B0 (n_6147), .Y
       (current_pc[6]));
  OAI2BB1X1 g89852__1881(.A0N (n_5997), .A1N (n_196), .B0 (n_6087), .Y
       (current_pc[18]));
  OAI2BB1X1 g89853__5115(.A0N (n_5997), .A1N (n_190), .B0 (n_6146), .Y
       (current_pc[15]));
  NAND4XL g89854__7482(.A (n_5617), .B (n_6034), .C (n_10531), .D
       (n_6161), .Y (n_6260));
  OAI2BB1X1 g89856__4733(.A0N (\genblk2.pcpi_div_quotient [17]), .A1N
       (n_5694), .B0 (n_6178), .Y (n_6259));
  OAI2BB1X1 g89857__6161(.A0N (\genblk2.pcpi_div_quotient [1]), .A1N
       (n_5694), .B0 (n_6193), .Y (n_6258));
  OAI2BB1X1 g89858__9315(.A0N (\genblk2.pcpi_div_dividend [2]), .A1N
       (n_5974), .B0 (n_6192), .Y (n_6257));
  OAI2BB1X1 g89859__9945(.A0N (\genblk2.pcpi_div_dividend [3]), .A1N
       (n_5974), .B0 (n_6191), .Y (n_6256));
  OAI2BB1X1 g89860__2883(.A0N (\genblk2.pcpi_div_dividend [4]), .A1N
       (n_5974), .B0 (n_6190), .Y (n_6255));
  OAI2BB1X1 g89861__2346(.A0N (\genblk2.pcpi_div_dividend [5]), .A1N
       (n_5974), .B0 (n_6189), .Y (n_6254));
  OAI2BB1X1 g89862__1666(.A0N (\genblk2.pcpi_div_dividend [6]), .A1N
       (n_5974), .B0 (n_6188), .Y (n_6253));
  OAI2BB1X1 g89863__7410(.A0N (\genblk2.pcpi_div_dividend [7]), .A1N
       (n_5974), .B0 (n_6187), .Y (n_6252));
  OAI2BB1X1 g89864__6417(.A0N (\genblk2.pcpi_div_quotient [8]), .A1N
       (n_5694), .B0 (n_6186), .Y (n_6251));
  OAI2BB1X1 g89865__5477(.A0N (\genblk2.pcpi_div_quotient [9]), .A1N
       (n_5694), .B0 (n_6185), .Y (n_6250));
  OAI2BB1X1 g89866__2398(.A0N (\genblk2.pcpi_div_quotient [10]), .A1N
       (n_5694), .B0 (n_6184), .Y (n_6249));
  OAI2BB1X1 g89867__5107(.A0N (\genblk2.pcpi_div_quotient [11]), .A1N
       (n_5694), .B0 (n_6183), .Y (n_6248));
  OAI2BB1X1 g89868__6260(.A0N (\genblk2.pcpi_div_quotient [12]), .A1N
       (n_5694), .B0 (n_6182), .Y (n_6247));
  OAI2BB1X1 g89869__4319(.A0N (\genblk2.pcpi_div_quotient [13]), .A1N
       (n_5694), .B0 (n_6181), .Y (n_6246));
  OAI2BB1X1 g89870__8428(.A0N (\genblk2.pcpi_div_quotient [14]), .A1N
       (n_5694), .B0 (n_6208), .Y (n_6245));
  OAI2BB1X1 g89871__5526(.A0N (\genblk2.pcpi_div_dividend [16]), .A1N
       (n_5974), .B0 (n_6195), .Y (n_6244));
  OAI2BB1X1 g89872__6783(.A0N (\genblk2.pcpi_div_quotient [18]), .A1N
       (n_5694), .B0 (n_6177), .Y (n_6243));
  OAI2BB1X1 g89873__3680(.A0N (\genblk2.pcpi_div_quotient [19]), .A1N
       (n_5694), .B0 (n_6176), .Y (n_6242));
  OAI2BB1X1 g89874__1617(.A0N (\genblk2.pcpi_div_quotient [20]), .A1N
       (n_5694), .B0 (n_6175), .Y (n_6241));
  OAI2BB1X1 g89875__2802(.A0N (\genblk2.pcpi_div_quotient [21]), .A1N
       (n_5694), .B0 (n_6165), .Y (n_6240));
  OAI2BB1X1 g89876__1705(.A0N (\genblk2.pcpi_div_quotient [22]), .A1N
       (n_5694), .B0 (n_6162), .Y (n_6239));
  OAI2BB1X1 g89877__5122(.A0N (\genblk2.pcpi_div_quotient [24]), .A1N
       (n_5694), .B0 (n_6196), .Y (n_6238));
  OAI2BB1X1 g89878__8246(.A0N (\genblk2.pcpi_div_quotient [25]), .A1N
       (n_5694), .B0 (n_6172), .Y (n_6237));
  OAI2BB1X1 g89879__7098(.A0N (\genblk2.pcpi_div_quotient [26]), .A1N
       (n_5694), .B0 (n_6171), .Y (n_6236));
  OAI2BB1X1 g89880__6131(.A0N (\genblk2.pcpi_div_quotient [27]), .A1N
       (n_5694), .B0 (n_6170), .Y (n_6235));
  OAI2BB1X1 g89881__1881(.A0N (\genblk2.pcpi_div_quotient [28]), .A1N
       (n_5694), .B0 (n_6169), .Y (n_6234));
  OAI2BB1X1 g89882__5115(.A0N (\genblk2.pcpi_div_quotient [29]), .A1N
       (n_5694), .B0 (n_6168), .Y (n_6233));
  OAI2BB1X1 g89883__7482(.A0N (\genblk2.pcpi_div_quotient [30]), .A1N
       (n_5694), .B0 (n_6167), .Y (n_6232));
  OAI2BB1X1 g89884__4733(.A0N (\genblk2.pcpi_div_quotient [31]), .A1N
       (n_5694), .B0 (n_6166), .Y (n_6231));
  OAI2BB1X1 g89885__6161(.A0N (\genblk2.pcpi_div_quotient [23]), .A1N
       (n_5694), .B0 (n_6173), .Y (n_6230));
  AOI22XL g89886__9315(.A0 (n_657), .A1 (mem_rdata[8]), .B0 (n_5998),
       .B1 (mem_rdata[24]), .Y (n_6229));
  MX2X1 g89887__9945(.A (reg_next_pc[1]), .B (n_160), .S0 (n_5997), .Y
       (current_pc[1]));
  NOR4X1 g89888__2883(.A (instr_beq), .B (instr_slli), .C (n_6064), .D
       (n_6127), .Y (n_6228));
  OR2X1 g89898__1666(.A (n_6532), .B (n_544), .Y (n_60));
  OAI2BB1X1 g89899__7410(.A0N (reg_out[2]), .A1N (n_5997), .B0
       (n_6152), .Y (n_6833));
  NOR2X1 g89901__5477(.A (n_5597), .B (n_6096), .Y (n_6224));
  NOR2BX1 g89902__2398(.AN (n_5597), .B (n_6096), .Y (n_6223));
  OAI2BB1X1 g89903__5107(.A0N (reg_out[3]), .A1N (n_5997), .B0
       (n_6151), .Y (n_6834));
  NAND2X1 g89904__6260(.A (n_228), .B (n_331), .Y (n_6222));
  OAI2BB1X1 g89905__4319(.A0N (reg_out[4]), .A1N (n_5997), .B0
       (n_6150), .Y (n_6835));
  NAND2X1 g89907__5526(.A (n_279), .B (n_6657), .Y (n_6220));
  NAND2X1 g89908__6783(.A (n_279), .B (n_6658), .Y (n_6219));
  NAND2X1 g89909__3680(.A (n_279), .B (n_6659), .Y (n_6218));
  NAND2X1 g89910__1617(.A (n_279), .B (n_6660), .Y (n_6217));
  NAND2X1 g89911__2802(.A (n_279), .B (n_6663), .Y (n_6216));
  NAND2X1 g89912__1705(.A (n_279), .B (n_6665), .Y (n_6215));
  NAND2X1 g89913__5122(.A (n_279), .B (n_6666), .Y (n_6214));
  NAND2X1 g89914__8246(.A (n_279), .B (n_6667), .Y (n_6213));
  NAND2X1 g89915__7098(.A (n_279), .B (n_6671), .Y (n_6212));
  NAND2X1 g89916__6131(.A (n_279), .B (n_6674), .Y (n_6211));
  OAI2BB1X1 g89917__1881(.A0N (reg_out[12]), .A1N (n_5997), .B0
       (n_6136), .Y (n_6843));
  OAI2BB1X1 g89918__5115(.A0N (reg_out[31]), .A1N (n_5997), .B0
       (n_6145), .Y (n_6862));
  OAI2BB1X1 g89919__7482(.A0N (reg_out[30]), .A1N (n_5997), .B0
       (n_6138), .Y (n_6861));
  OAI2BB1X1 g89920__4733(.A0N (reg_out[29]), .A1N (n_5997), .B0
       (n_6135), .Y (n_6860));
  OAI2BB1X1 g89921__6161(.A0N (reg_out[28]), .A1N (n_5997), .B0
       (n_6148), .Y (n_6859));
  OAI2BB1X1 g89922__9315(.A0N (reg_out[27]), .A1N (n_5997), .B0
       (n_6133), .Y (n_6858));
  OAI2BB1X1 g89923__9945(.A0N (reg_out[26]), .A1N (n_5997), .B0
       (n_6131), .Y (n_6857));
  OAI2BB1X1 g89924__2883(.A0N (reg_out[25]), .A1N (n_5997), .B0
       (n_6129), .Y (n_6856));
  OAI2BB1X1 g89925__2346(.A0N (reg_out[24]), .A1N (n_5997), .B0
       (n_6128), .Y (n_6855));
  OAI2BB1X1 g89926__1666(.A0N (reg_out[23]), .A1N (n_5997), .B0
       (n_6100), .Y (n_6854));
  OAI2BB1X1 g89927__7410(.A0N (reg_out[22]), .A1N (n_5997), .B0
       (n_6093), .Y (n_6853));
  OAI2BB1X1 g89928__6417(.A0N (reg_out[21]), .A1N (n_5997), .B0
       (n_6102), .Y (n_6852));
  OAI2BB1X1 g89929__5477(.A0N (reg_out[20]), .A1N (n_5997), .B0
       (n_6099), .Y (n_6851));
  OAI2BB1X1 g89930__2398(.A0N (reg_out[19]), .A1N (n_5997), .B0
       (n_6089), .Y (n_6850));
  OAI2BB1X1 g89931__5107(.A0N (reg_out[18]), .A1N (n_5997), .B0
       (n_6087), .Y (n_6849));
  OAI2BB1X1 g89932__6260(.A0N (reg_out[17]), .A1N (n_5997), .B0
       (n_6084), .Y (n_6848));
  OAI2BB1X1 g89933__4319(.A0N (reg_out[16]), .A1N (n_5997), .B0
       (n_6083), .Y (n_6847));
  OAI2BB1X1 g89934__8428(.A0N (reg_out[15]), .A1N (n_5997), .B0
       (n_6146), .Y (n_6846));
  OAI2BB1X1 g89935__5526(.A0N (reg_out[14]), .A1N (n_5997), .B0
       (n_6130), .Y (n_6845));
  OAI2BB1X1 g89936__6783(.A0N (reg_out[13]), .A1N (n_5997), .B0
       (n_6132), .Y (n_6844));
  OAI2BB1X1 g89937__3680(.A0N (reg_out[11]), .A1N (n_5997), .B0
       (n_6137), .Y (n_6842));
  OAI2BB1X1 g89938__1617(.A0N (reg_out[10]), .A1N (n_5997), .B0
       (n_6140), .Y (n_6841));
  OAI2BB1X1 g89939__2802(.A0N (reg_out[9]), .A1N (n_5997), .B0
       (n_6142), .Y (n_6840));
  OAI2BB1X1 g89940__1705(.A0N (reg_out[8]), .A1N (n_5997), .B0
       (n_6143), .Y (n_6839));
  OAI2BB1X1 g89942__8246(.A0N (reg_out[7]), .A1N (n_5997), .B0
       (n_6144), .Y (n_6838));
  OAI2BB1X1 g89943__7098(.A0N (reg_out[6]), .A1N (n_5997), .B0
       (n_6147), .Y (n_6837));
  OAI2BB1X1 g89944__6131(.A0N (reg_out[5]), .A1N (n_5997), .B0
       (n_6149), .Y (n_6836));
  OR2X1 g89945__1881(.A (pcpi_timeout_counter[3]), .B (n_218), .Y
       (n_258));
  NOR4X1 g89946__5115(.A (instr_add), .B (instr_addi), .C (n_6029), .D
       (n_6085), .Y (n_6227));
  NAND2BX1 g89947__7482(.AN (n_6050), .B (n_6554), .Y (n_158));
  AOI22XL g89949__4733(.A0 (\genblk2.pcpi_div_dividend [14]), .A1
       (n_5974), .B0 (\genblk2.pcpi_div_outsign ), .B1
       (\genblk2.pcpi_div_n_2159 ), .Y (n_6208));
  OAI2BB1X1 g89956__7410(.A0N (n_6058), .A1N (n_6052), .B0 (resetn), .Y
       (n_6201));
  AOI22XL g89961__6260(.A0 (\genblk2.pcpi_div_dividend [24]), .A1
       (n_5974), .B0 (\genblk2.pcpi_div_outsign ), .B1
       (\genblk2.pcpi_div_n_2149 ), .Y (n_6196));
  AOI22XL g89962__4319(.A0 (\genblk2.pcpi_div_quotient [16]), .A1
       (n_5694), .B0 (\genblk2.pcpi_div_outsign ), .B1
       (\genblk2.pcpi_div_n_2157 ), .Y (n_6195));
  AOI22XL g89964__5526(.A0 (\genblk2.pcpi_div_dividend [1]), .A1
       (n_5974), .B0 (\genblk2.pcpi_div_outsign ), .B1
       (\genblk2.pcpi_div_n_2172 ), .Y (n_6193));
  AOI22XL g89965__6783(.A0 (\genblk2.pcpi_div_quotient [2]), .A1
       (n_5694), .B0 (\genblk2.pcpi_div_outsign ), .B1
       (\genblk2.pcpi_div_n_2171 ), .Y (n_6192));
  AOI22XL g89966__3680(.A0 (\genblk2.pcpi_div_quotient [3]), .A1
       (n_5694), .B0 (\genblk2.pcpi_div_outsign ), .B1
       (\genblk2.pcpi_div_n_2170 ), .Y (n_6191));
  AOI22XL g89967__1617(.A0 (\genblk2.pcpi_div_quotient [4]), .A1
       (n_5694), .B0 (\genblk2.pcpi_div_outsign ), .B1
       (\genblk2.pcpi_div_n_2169 ), .Y (n_6190));
  AOI22XL g89968__2802(.A0 (\genblk2.pcpi_div_quotient [5]), .A1
       (n_5694), .B0 (\genblk2.pcpi_div_outsign ), .B1
       (\genblk2.pcpi_div_n_2168 ), .Y (n_6189));
  AOI22XL g89969__1705(.A0 (\genblk2.pcpi_div_quotient [6]), .A1
       (n_5694), .B0 (\genblk2.pcpi_div_outsign ), .B1
       (\genblk2.pcpi_div_n_2167 ), .Y (n_6188));
  AOI22XL g89970__5122(.A0 (\genblk2.pcpi_div_quotient [7]), .A1
       (n_5694), .B0 (\genblk2.pcpi_div_outsign ), .B1
       (\genblk2.pcpi_div_n_2166 ), .Y (n_6187));
  AOI22XL g89971__8246(.A0 (\genblk2.pcpi_div_dividend [8]), .A1
       (n_5974), .B0 (\genblk2.pcpi_div_outsign ), .B1
       (\genblk2.pcpi_div_n_2165 ), .Y (n_6186));
  AOI22XL g89972__7098(.A0 (\genblk2.pcpi_div_dividend [9]), .A1
       (n_5974), .B0 (\genblk2.pcpi_div_outsign ), .B1
       (\genblk2.pcpi_div_n_2164 ), .Y (n_6185));
  AOI22XL g89973__6131(.A0 (\genblk2.pcpi_div_dividend [10]), .A1
       (n_5974), .B0 (\genblk2.pcpi_div_outsign ), .B1
       (\genblk2.pcpi_div_n_2163 ), .Y (n_6184));
  AOI22XL g89974__1881(.A0 (\genblk2.pcpi_div_dividend [11]), .A1
       (n_5974), .B0 (\genblk2.pcpi_div_outsign ), .B1
       (\genblk2.pcpi_div_n_2162 ), .Y (n_6183));
  AOI22XL g89975__5115(.A0 (\genblk2.pcpi_div_dividend [12]), .A1
       (n_5974), .B0 (\genblk2.pcpi_div_outsign ), .B1
       (\genblk2.pcpi_div_n_2161 ), .Y (n_6182));
  AOI22XL g89976__7482(.A0 (\genblk2.pcpi_div_dividend [13]), .A1
       (n_5974), .B0 (\genblk2.pcpi_div_outsign ), .B1
       (\genblk2.pcpi_div_n_2160 ), .Y (n_6181));
  AOI22XL g89978__6161(.A0 (\genblk2.pcpi_div_dividend [15]), .A1
       (n_5974), .B0 (\genblk2.pcpi_div_outsign ), .B1
       (\genblk2.pcpi_div_n_2158 ), .Y (n_6179));
  AOI22XL g89979__9315(.A0 (\genblk2.pcpi_div_dividend [17]), .A1
       (n_5974), .B0 (\genblk2.pcpi_div_outsign ), .B1
       (\genblk2.pcpi_div_n_2156 ), .Y (n_6178));
  AOI22XL g89980__9945(.A0 (\genblk2.pcpi_div_dividend [18]), .A1
       (n_5974), .B0 (\genblk2.pcpi_div_outsign ), .B1
       (\genblk2.pcpi_div_n_2155 ), .Y (n_6177));
  AOI22XL g89981__2883(.A0 (\genblk2.pcpi_div_dividend [19]), .A1
       (n_5974), .B0 (\genblk2.pcpi_div_outsign ), .B1
       (\genblk2.pcpi_div_n_2154 ), .Y (n_6176));
  AOI22XL g89982__2346(.A0 (\genblk2.pcpi_div_dividend [20]), .A1
       (n_5974), .B0 (\genblk2.pcpi_div_outsign ), .B1
       (\genblk2.pcpi_div_n_2153 ), .Y (n_6175));
  AOI22XL g89984__7410(.A0 (\genblk2.pcpi_div_dividend [23]), .A1
       (n_5974), .B0 (\genblk2.pcpi_div_outsign ), .B1
       (\genblk2.pcpi_div_n_2150 ), .Y (n_6173));
  AOI22XL g89985__6417(.A0 (\genblk2.pcpi_div_dividend [25]), .A1
       (n_5974), .B0 (\genblk2.pcpi_div_outsign ), .B1
       (\genblk2.pcpi_div_n_2148 ), .Y (n_6172));
  AOI22XL g89986__5477(.A0 (\genblk2.pcpi_div_dividend [26]), .A1
       (n_5974), .B0 (\genblk2.pcpi_div_outsign ), .B1
       (\genblk2.pcpi_div_n_2147 ), .Y (n_6171));
  AOI22XL g89987__2398(.A0 (\genblk2.pcpi_div_dividend [27]), .A1
       (n_5974), .B0 (\genblk2.pcpi_div_outsign ), .B1
       (\genblk2.pcpi_div_n_2146 ), .Y (n_6170));
  AOI22XL g89988__5107(.A0 (\genblk2.pcpi_div_dividend [28]), .A1
       (n_5974), .B0 (\genblk2.pcpi_div_outsign ), .B1
       (\genblk2.pcpi_div_n_2145 ), .Y (n_6169));
  AOI22XL g89989__6260(.A0 (\genblk2.pcpi_div_dividend [29]), .A1
       (n_5974), .B0 (\genblk2.pcpi_div_outsign ), .B1
       (\genblk2.pcpi_div_n_2144 ), .Y (n_6168));
  AOI22XL g89990__4319(.A0 (\genblk2.pcpi_div_dividend [30]), .A1
       (n_5974), .B0 (\genblk2.pcpi_div_outsign ), .B1
       (\genblk2.pcpi_div_n_2143 ), .Y (n_6167));
  AOI22XL g89991__8428(.A0 (\genblk2.pcpi_div_dividend [31]), .A1
       (n_5974), .B0 (\genblk2.pcpi_div_outsign ), .B1
       (\genblk2.pcpi_div_n_2142 ), .Y (n_6166));
  AOI22XL g89992__5526(.A0 (\genblk2.pcpi_div_dividend [21]), .A1
       (n_5974), .B0 (\genblk2.pcpi_div_outsign ), .B1
       (\genblk2.pcpi_div_n_2152 ), .Y (n_6165));
  AOI22XL g89995__1617(.A0 (\genblk2.pcpi_div_dividend [22]), .A1
       (n_5974), .B0 (\genblk2.pcpi_div_outsign ), .B1
       (\genblk2.pcpi_div_n_2151 ), .Y (n_6162));
  NOR4X1 g89996__2802(.A (n_5588), .B (n_5587), .C (n_6057), .D
       (n_10491), .Y (n_6161));
  OAI22X1 g89997__1705(.A0 (reg_out[1]), .A1 (n_320), .B0
       (reg_next_pc[1]), .B1 (n_5997), .Y (n_6160));
  OAI31X1 g90005__4733(.A0 (reg_op1[0]), .A1 (n_565), .A2 (n_5984), .B0
       (n_228), .Y (n_340));
  NOR2X1 g90007__6161(.A (n_577), .B (n_313), .Y (n_61756_BAR));
  NOR2BX1 g90011__2346(.AN (\reg_op2[1]_9670 ), .B (n_608), .Y
       (n_6124));
  NOR2X1 g90015__5477(.A (n_42), .B (n_5984), .Y (n_6122));
  NOR2X1 g90017__5107(.A (n_634), .B (n_313), .Y (n_61792_BAR));
  NOR2BX1 g90020__8428(.AN (\reg_op2[18]_9687 ), .B (n_6517), .Y
       (n_6121));
  NOR2X1 g90025__2802(.A (n_5829), .B (n_313), .Y (n_61806_BAR));
  NOR2X1 g90026__1705(.A (n_5786), .B (n_313), .Y (n_61804_BAR));
  NOR2X1 g90028__8246(.A (n_5827), .B (n_313), .Y (n_61798_BAR));
  NOR2BX1 g90030__6131(.AN (\reg_op2[7]_9676 ), .B (n_608), .Y
       (n_6119));
  NOR2X1 g90034__4733(.A (n_5813), .B (n_313), .Y (n_61784_BAR));
  NOR2X1 g90042__6417(.A (n_5859), .B (n_313), .Y (n_61762_BAR));
  NOR2BX1 g90043__5477(.AN (\reg_op2[23]_9692 ), .B (n_6517), .Y
       (n_6118));
  NOR2X1 g90044__2398(.A (n_717), .B (n_313), .Y (n_61760_BAR));
  NOR2X1 g90045__5107(.A (n_578), .B (n_313), .Y (n_61758_BAR));
  NOR2BX1 g90046__6260(.AN (\reg_op2[19]_9688 ), .B (n_6517), .Y
       (n_6117));
  NOR2BX1 g90048__8428(.AN (\reg_op2[0]_9669 ), .B (n_608), .Y
       (n_6115));
  NOR2BX1 g90049__5526(.AN (\reg_op2[6]_9675 ), .B (n_608), .Y
       (n_6114));
  NOR2BX1 g90050__6783(.AN (\reg_op2[16]_9685 ), .B (n_6517), .Y
       (n_6113));
  NOR2BX1 g90051__3680(.AN (\reg_op2[22]_9691 ), .B (n_6517), .Y
       (n_6112));
  NOR2BX1 g90052__1617(.AN (\reg_op2[17]_9686 ), .B (n_6517), .Y
       (n_6111));
  NOR2BX1 g90053__2802(.AN (\reg_op2[20]_9689 ), .B (n_6517), .Y
       (n_6110));
  NOR2BX1 g90057__7098(.AN (\reg_op2[21]_9690 ), .B (n_6517), .Y
       (n_6106));
  NAND2XL g90058__6131(.A (reg_next_pc[2]), .B (n_320), .Y (n_6152));
  NAND2XL g90059__1881(.A (reg_next_pc[3]), .B (n_320), .Y (n_6151));
  NAND2XL g90060__5115(.A (reg_next_pc[4]), .B (n_320), .Y (n_6150));
  NAND2XL g90061__7482(.A (reg_next_pc[5]), .B (n_320), .Y (n_6149));
  NAND2XL g90062__4733(.A (reg_next_pc[28]), .B (n_320), .Y (n_6148));
  NAND2XL g90063__6161(.A (reg_next_pc[6]), .B (n_320), .Y (n_6147));
  NAND2BXL g90064__9315(.AN (n_222), .B (prefetched_high_word), .Y
       (n_6531));
  NAND2XL g90065__9945(.A (reg_next_pc[15]), .B (n_320), .Y (n_6146));
  NAND2XL g90066__2883(.A (reg_next_pc[31]), .B (n_320), .Y (n_6145));
  NAND2XL g90067__2346(.A (reg_next_pc[7]), .B (n_320), .Y (n_6144));
  NAND2XL g90068__1666(.A (reg_next_pc[8]), .B (n_320), .Y (n_6143));
  NAND2XL g90069__7410(.A (reg_next_pc[9]), .B (n_320), .Y (n_6142));
  NOR2BX1 g90070__6417(.AN (\reg_op2[6]_9675 ), .B (n_5984), .Y
       (n_6141));
  NAND2XL g90071__5477(.A (reg_next_pc[10]), .B (n_320), .Y (n_6140));
  NAND2XL g90073__5107(.A (reg_next_pc[30]), .B (n_320), .Y (n_6138));
  NAND2XL g90074__6260(.A (reg_next_pc[11]), .B (n_320), .Y (n_6137));
  NAND2XL g90075__4319(.A (reg_next_pc[12]), .B (n_320), .Y (n_6136));
  NAND2XL g90076__8428(.A (reg_next_pc[29]), .B (n_320), .Y (n_6135));
  NOR2BX1 g90077__5526(.AN (\reg_op2[0]_9669 ), .B (n_5984), .Y
       (n_6134));
  NAND2XL g90078__6783(.A (reg_next_pc[27]), .B (n_320), .Y (n_6133));
  NAND2XL g90079__3680(.A (reg_next_pc[13]), .B (n_320), .Y (n_6132));
  NAND2XL g90080__1617(.A (reg_next_pc[26]), .B (n_320), .Y (n_6131));
  NAND2XL g90081__2802(.A (reg_next_pc[14]), .B (n_320), .Y (n_6130));
  NAND2XL g90082__1705(.A (reg_next_pc[25]), .B (n_320), .Y (n_6129));
  NAND2XL g90083__5122(.A (reg_next_pc[24]), .B (n_320), .Y (n_6128));
  NAND2BX1 g90084__8246(.AN (instr_bltu), .B (n_6058), .Y (n_6127));
  INVX1 g90085(.A (n_6094), .Y (n_6095));
  INVX1 g90086(.A (n_6082), .Y (n_122));
  INVX1 g90087(.A (n_311), .Y (n_657));
  NOR2X1 g90096__9315(.A (n_756), .B (n_608), .Y (n_6073));
  NOR2X1 g90097__9945(.A (\genblk2.pcpi_div_minus_2470_59_n_477 ), .B
       (n_608), .Y (n_6072));
  NOR2X1 g90098__2883(.A (n_725), .B (n_608), .Y (n_6071));
  NOR2X1 g90099__2346(.A (\genblk2.pcpi_div_minus_2470_59_n_487 ), .B
       (n_608), .Y (n_6070));
  NOR3BX1 g90101__7410(.AN (mem_valid_9465), .B (mem_ready), .C
       (n_544), .Y (n_6068));
  OAI21X1 g90102__6417(.A0 (compressed_instr), .A1 (instr_jal), .B0
       (n_6045), .Y (n_6606));
  AOI22XL g90103__5477(.A0 (count_instr[0]), .A1 (instr_rdinstr), .B0
       (instr_rdinstrh), .B1 (count_instr[32]), .Y (n_6067));
  AOI22XL g90104__2398(.A0 (count_cycle[0]), .A1 (instr_rdcycle), .B0
       (instr_rdcycleh), .B1 (count_cycle[32]), .Y (n_6066));
  MX2X1 g90106__6260(.A (compressed_instr), .B (decoded_imm_j[1]), .S0
       (instr_jal), .Y (n_6605));
  OR4X1 g90107__4319(.A (instr_srl), .B (instr_sra), .C (instr_bge), .D
       (instr_bne), .Y (n_6064));
  XNOR2X1 g90108__8428(.A (cpu_state[1]), .B (cpu_state[0]), .Y
       (n_6063));
  NOR4X1 g90110__6783(.A (instr_srli), .B (instr_srai), .C (instr_sb),
       .D (instr_lb), .Y (n_6061));
  NOR2BX1 g90111__3680(.AN (\reg_op2[7]_9676 ), .B (n_5984), .Y
       (n_6105));
  XNOR2X1 g90112__1617(.A (\reg_op2[16]_9685 ), .B (n_5813), .Y
       (n_6661));
  NOR2X1 g90113__2802(.A (\genblk2.pcpi_div_minus_2470_59_n_477 ), .B
       (n_5984), .Y (n_6104));
  NOR2X1 g90114__1705(.A (\genblk2.pcpi_div_minus_2470_59_n_487 ), .B
       (n_5984), .Y (n_6103));
  OR2X1 g90115__5122(.A (pcpi_timeout_counter[2]), .B (n_162), .Y
       (n_218));
  NAND2XL g90116__8246(.A (reg_next_pc[21]), .B (n_320), .Y (n_6102));
  NOR2X1 g90117__7098(.A (n_725), .B (n_5984), .Y (n_6101));
  NAND2XL g90118__6131(.A (reg_next_pc[23]), .B (n_320), .Y (n_6100));
  NAND2XL g90119__1881(.A (reg_next_pc[20]), .B (n_320), .Y (n_6099));
  NOR2X1 g90120__5115(.A (n_756), .B (n_5984), .Y (n_6098));
  XNOR2X1 g90121__7482(.A (\reg_op2[24]_9693 ), .B (n_713), .Y
       (n_6668));
  NAND2X1 g90122__4733(.A (n_6552), .B (n_6553), .Y (n_6674));
  NAND2X1 g90123__6161(.A (n_6550), .B (n_6551), .Y (n_6671));
  NAND2X1 g90124__9315(.A (n_138), .B (n_6546), .Y (n_6667));
  NAND2X1 g90125__9945(.A (n_6547), .B (n_6544), .Y (n_6666));
  NAND2X1 g90126__2883(.A (n_152), .B (n_6543), .Y (n_6665));
  NAND2X1 g90127__2346(.A (n_136), .B (n_6548), .Y (n_6663));
  NOR2BX1 g90128__1666(.AN (\reg_op2[1]_9670 ), .B (n_5984), .Y
       (n_6097));
  NAND2X1 g90129__7410(.A (n_6534), .B (n_6538), .Y (n_6659));
  NAND2X1 g90130__6417(.A (n_6535), .B (n_6559), .Y (n_6658));
  NAND3BXL g90131__5477(.AN (n_6530), .B (n_5599), .C (n_5598), .Y
       (n_6096));
  NAND2X1 g90132__2398(.A (n_6533), .B (n_6537), .Y (n_6657));
  NAND3X1 g90133__5107(.A (mem_do_rinst), .B (mem_state[1]), .C
       (mem_state[0]), .Y (n_6567));
  XNOR2X1 g90134__6260(.A (\reg_op2[28]_9697 ), .B (n_5788), .Y
       (n_6672));
  NOR3X1 g90135__4319(.A (instr_lw), .B (instr_lhu), .C (instr_lbu), .Y
       (n_6094));
  NAND2XL g90136__8428(.A (reg_next_pc[22]), .B (n_320), .Y (n_6093));
  XNOR2X1 g90137__5526(.A (\reg_op2[29]_9698 ), .B (n_716), .Y
       (n_6673));
  OA21X1 g90138__6783(.A0 (\reg_op2[26]_9695 ), .A1 (n_5786), .B0
       (n_6549), .Y (n_6092));
  OA21X1 g90139__3680(.A0 (\reg_op2[25]_9694 ), .A1 (n_5784), .B0
       (n_156), .Y (n_6091));
  OA21X1 g90140__1617(.A0 (\reg_op2[20]_9689 ), .A1 (n_634), .B0
       (n_6542), .Y (n_6090));
  NAND2XL g90141__2802(.A (reg_next_pc[19]), .B (n_320), .Y (n_6089));
  OA21X1 g90142__1705(.A0 (\reg_op2[17]_9686 ), .A1 (n_715), .B0
       (n_154), .Y (n_6088));
  NAND2X1 g90143__5122(.A (n_6536), .B (n_6541), .Y (n_6660));
  NAND2BX1 g90144__8246(.AN (n_6050), .B (mem_do_wdata), .Y (n_6532));
  OR2X1 g90145__7098(.A (mem_do_rdata), .B (n_313), .Y (n_6554));
  MX2X1 g90146__6131(.A (reg_out[15]), .B (alu_out_q[15]), .S0
       (latched_stalu), .Y (n_190));
  MX2X1 g90147__1881(.A (reg_out[14]), .B (alu_out_q[14]), .S0
       (latched_stalu), .Y (n_188));
  MX2X1 g90148__5115(.A (reg_out[13]), .B (alu_out_q[13]), .S0
       (latched_stalu), .Y (n_172));
  MX2X1 g90149__7482(.A (reg_out[12]), .B (alu_out_q[12]), .S0
       (latched_stalu), .Y (n_186));
  MX2X1 g90150__4733(.A (reg_out[11]), .B (alu_out_q[11]), .S0
       (latched_stalu), .Y (n_184));
  MX2X1 g90151__6161(.A (reg_out[10]), .B (alu_out_q[10]), .S0
       (latched_stalu), .Y (n_182));
  MX2X1 g90152__9315(.A (reg_out[9]), .B (alu_out_q[9]), .S0
       (latched_stalu), .Y (n_180));
  MX2X1 g90153__9945(.A (reg_out[7]), .B (alu_out_q[7]), .S0
       (latched_stalu), .Y (n_176));
  MX2X1 g90154__2883(.A (reg_out[6]), .B (alu_out_q[6]), .S0
       (latched_stalu), .Y (n_174));
  MX2X1 g90155__2346(.A (reg_out[1]), .B (alu_out_q[1]), .S0
       (latched_stalu), .Y (n_160));
  MX2X1 g90156__1666(.A (reg_out[8]), .B (alu_out_q[8]), .S0
       (latched_stalu), .Y (n_178));
  MX2X1 g90157__7410(.A (reg_out[18]), .B (alu_out_q[18]), .S0
       (latched_stalu), .Y (n_196));
  NAND2XL g90158__6417(.A (reg_next_pc[18]), .B (n_320), .Y (n_6087));
  NAND2BX1 g90159__5477(.AN (instr_blt), .B (n_6052), .Y (n_6086));
  OR2X1 g90160__2398(.A (instr_jal), .B (n_6514), .Y (n_6085));
  NAND2XL g90161__5107(.A (reg_next_pc[17]), .B (n_320), .Y (n_6084));
  NAND2XL g90162__6260(.A (reg_next_pc[16]), .B (n_320), .Y (n_6083));
  NAND2X1 g90163__4319(.A (\reg_op1[1]_9638 ), .B (n_5980), .Y (n_228));
  AOI21X1 g90164__8428(.A0 (mem_wordsize[0]), .A1 (\reg_op1[1]_9638 ),
       .B0 (mem_wordsize[1]), .Y (n_6082));
  NAND3X1 g90165__5526(.A (reg_op1[0]), .B (n_565), .C (n_5996), .Y
       (n_311));
  NAND3X1 g90166__6783(.A (\reg_op1[1]_9638 ), .B (reg_op1[0]), .C
       (n_5996), .Y (n_331));
  NAND2X1 g90234__3680(.A (n_5586), .B (n_5585), .Y (n_6057));
  NOR2X1 g90235__1617(.A (\reg_op1[17]_9654 ), .B (\reg_op2[17]_9686 ),
       .Y (n_6056));
  NOR2X1 g90236__2802(.A (\reg_op1[5]_9642 ), .B (\reg_op2[5]_9674 ),
       .Y (n_6055));
  NOR2X1 g90237__1705(.A (\reg_op1[22]_9659 ), .B (\reg_op2[22]_9691 ),
       .Y (n_6054));
  OR2X1 g90238__5122(.A (cpu_state[3]), .B (cpu_state[5]), .Y
       (n_14409_BAR));
  NOR2X1 g90239__8246(.A (\reg_op1[16]_9653 ), .B (\reg_op2[16]_9685 ),
       .Y (n_6053));
  NAND2X1 g90240__7098(.A (mem_valid_9465), .B (mem_ready), .Y
       (n_6060));
  NAND2X1 g90241__6131(.A (\reg_op2[31]_9700 ), .B (\reg_op1[31]_9668
       ), .Y (n_6059));
  NAND2X1 g90242__1881(.A (n_628), .B (n_565), .Y (n_42));
  NOR2XL g90243__5115(.A (instr_sltu), .B (instr_sltiu), .Y (n_6058));
  OR2X2 g90244__7482(.A (n_6026), .B (n_555), .Y (n_320));
  INVX2 g90247(.A (n_6048), .Y (n_283));
  NAND2XL g90251__4733(.A (decoded_imm_j[2]), .B (instr_jal), .Y
       (n_6045));
  NOR2X1 g90252__6161(.A (\reg_op1[29]_9666 ), .B (\reg_op2[29]_9698 ),
       .Y (n_6044));
  NOR2X1 g90253__9315(.A (\reg_op1[28]_9665 ), .B (\reg_op2[28]_9697 ),
       .Y (n_6043));
  NOR2XL g90254__9945(.A (instr_sll), .B (instr_lh), .Y (n_6042));
  AND2X1 g90255__2883(.A (decoded_imm_j[20]), .B (instr_jal), .Y
       (n_6624));
  AND2X1 g90256__2346(.A (instr_jal), .B (decoded_imm_j[19]), .Y
       (n_6623));
  AND2X1 g90257__1666(.A (instr_jal), .B (decoded_imm_j[18]), .Y
       (n_6622));
  AND2X1 g90258__7410(.A (instr_jal), .B (decoded_imm_j[17]), .Y
       (n_6621));
  AND2X1 g90259__6417(.A (instr_jal), .B (decoded_imm_j[16]), .Y
       (n_6620));
  AND2X1 g90260__5477(.A (instr_jal), .B (decoded_imm_j[15]), .Y
       (n_6619));
  AND2X1 g90261__2398(.A (instr_jal), .B (decoded_imm_j[14]), .Y
       (n_6618));
  AND2X1 g90262__5107(.A (instr_jal), .B (decoded_imm_j[13]), .Y
       (n_6617));
  AND2X1 g90263__6260(.A (instr_jal), .B (decoded_imm_j[12]), .Y
       (n_6616));
  AND2X1 g90264__4319(.A (instr_jal), .B (decoded_imm_j[11]), .Y
       (n_6615));
  AND2X1 g90265__8428(.A (instr_jal), .B (decoded_imm_j[10]), .Y
       (n_6614));
  NOR2X1 g90266__5526(.A (\reg_op1[27]_9664 ), .B (\reg_op2[27]_9696 ),
       .Y (n_6041));
  AND2X1 g90267__6783(.A (instr_jal), .B (decoded_imm_j[4]), .Y
       (n_6608));
  AND2X1 g90268__3680(.A (instr_jal), .B (decoded_imm_j[3]), .Y
       (n_6607));
  NOR2X1 g90269__1617(.A (\reg_op1[19]_9656 ), .B (\reg_op2[19]_9688 ),
       .Y (n_6040));
  AND2X1 g90270__2802(.A (instr_jal), .B (decoded_imm_j[5]), .Y
       (n_6609));
  NOR2X1 g90271__1705(.A (\reg_op1[21]_9658 ), .B (\reg_op2[21]_9690 ),
       .Y (n_6039));
  NOR2X1 g90272__5122(.A (\reg_op1[25]_9662 ), .B (\reg_op2[25]_9694 ),
       .Y (n_6038));
  NOR2X1 g90273__8246(.A (\reg_op1[3]_9640 ), .B (\reg_op2[3]_9672 ),
       .Y (n_6037));
  NOR2X1 g90274__7098(.A (\reg_op1[30]_9667 ), .B (\reg_op2[30]_9699 ),
       .Y (n_6036));
  AND2X1 g90275__6131(.A (instr_jal), .B (decoded_imm_j[8]), .Y
       (n_6612));
  AND2X1 g90276__1881(.A (instr_jal), .B (decoded_imm_j[6]), .Y
       (n_6610));
  NOR2X1 g90277__5115(.A (\reg_op1[2]_9639 ), .B (\reg_op2[2]_9671 ),
       .Y (n_6035));
  AND2X1 g90278__7482(.A (instr_jal), .B (decoded_imm_j[9]), .Y
       (n_6613));
  NOR2XL g90279__4733(.A (n_5616), .B (n_5615), .Y (n_6034));
  NOR2X1 g90280__6161(.A (\reg_op1[26]_9663 ), .B (\reg_op2[26]_9695 ),
       .Y (n_6033));
  NOR2X1 g90281__9315(.A (\reg_op1[24]_9661 ), .B (\reg_op2[24]_9693 ),
       .Y (n_6032));
  AND2X1 g90282__9945(.A (instr_jal), .B (decoded_imm_j[7]), .Y
       (n_6611));
  NOR2X1 g90283__2883(.A (\reg_op1[23]_9660 ), .B (\reg_op2[23]_9692 ),
       .Y (n_6031));
  NOR2X1 g90284__2346(.A (\reg_op1[20]_9657 ), .B (\reg_op2[20]_9689 ),
       .Y (n_6030));
  OR2X1 g90285__1666(.A (instr_jalr), .B (instr_sub), .Y (n_6029));
  NOR2X1 g90286__7410(.A (\reg_op1[4]_9641 ), .B (\reg_op2[4]_9673 ),
       .Y (n_6028));
  NAND2X1 g90287__6417(.A (\reg_op2[20]_9689 ), .B (n_634), .Y
       (n_6542));
  NAND2X1 g90288__5477(.A (\reg_op1[5]_9642 ), .B (n_756), .Y (n_6536));
  NAND2X1 g90289__2398(.A (\reg_op2[4]_9673 ), .B (n_717), .Y (n_6538));
  NAND2X1 g90290__5107(.A (\reg_op2[5]_9674 ), .B (n_5859), .Y
       (n_6541));
  NAND2X1 g90291__6260(.A (n_555), .B (resetn), .Y (n_222));
  NAND2X1 g90292__4319(.A (\reg_op1[3]_9640 ), .B (n_725), .Y (n_6535));
  NAND2X1 g90293__8428(.A (\reg_op2[30]_9699 ), .B (n_718), .Y
       (n_6552));
  NAND2X1 g90294__5526(.A (\reg_op2[23]_9692 ), .B (n_5827), .Y
       (n_138));
  NAND2BX1 g90295__6783(.AN (\reg_op2[23]_9692 ), .B (\reg_op1[23]_9660
       ), .Y (n_6546));
  NAND2BX1 g90296__3680(.AN (\reg_op2[22]_9691 ), .B (\reg_op1[22]_9659
       ), .Y (n_6544));
  NAND2X1 g90297__1617(.A (\reg_op2[21]_9690 ), .B (n_637), .Y (n_152));
  NAND2BX1 g90298__2802(.AN (\reg_op2[21]_9690 ), .B (\reg_op1[21]_9658
       ), .Y (n_6543));
  NAND2X1 g90299__1705(.A (\reg_op2[19]_9688 ), .B (n_747), .Y (n_136));
  NAND2BX1 g90300__5122(.AN (\reg_op2[19]_9688 ), .B (\reg_op1[19]_9656
       ), .Y (n_6548));
  OR2X1 g90301__8246(.A (mem_do_wdata), .B (mem_do_rdata), .Y (n_6555));
  OR2X1 g90302__7098(.A (pcpi_timeout_counter[0]), .B
       (pcpi_timeout_counter[1]), .Y (n_162));
  NAND2X1 g90303__6131(.A (\reg_op2[22]_9691 ), .B (n_576), .Y
       (n_6547));
  NAND2BX1 g90304__1881(.AN (\reg_op2[27]_9696 ), .B (\reg_op1[27]_9664
       ), .Y (n_6551));
  NAND2X1 g90305__5115(.A (\reg_op2[27]_9696 ), .B (n_5829), .Y
       (n_6550));
  NAND2X1 g90306__7482(.A (\reg_op2[26]_9695 ), .B (n_5786), .Y
       (n_6549));
  NAND2BX1 g90307__4733(.AN (\reg_op2[30]_9699 ), .B (\reg_op1[30]_9667
       ), .Y (n_6553));
  NAND2XL g90308__6161(.A (is_beq_bne_blt_bge_bltu_bgeu), .B (resetn),
       .Y (n_130));
  NAND2X1 g90309__9315(.A (\reg_op2[17]_9686 ), .B (n_715), .Y (n_154));
  NAND2X1 g90310__9945(.A (\reg_op1[4]_9641 ), .B
       (\genblk2.pcpi_div_minus_2470_59_n_477 ), .Y (n_6534));
  NOR2XL g90311__2883(.A (instr_slt), .B (instr_slti), .Y (n_6052));
  OR2X1 g90312__2346(.A (instr_auipc), .B (instr_lui), .Y (n_6514));
  NAND2X1 g90313__1666(.A (\reg_op2[3]_9672 ), .B (n_578), .Y (n_6559));
  NAND2X1 g90314__7410(.A (\reg_op2[25]_9694 ), .B (n_5784), .Y
       (n_156));
  NOR2X1 g90315__6417(.A (\reg_op1[31]_9668 ), .B (\reg_op2[31]_9700 ),
       .Y (n_6051));
  NAND2X1 g90316__5477(.A (\reg_op2[2]_9671 ), .B (n_577), .Y (n_6537));
  NAND2X1 g90317__2398(.A (\reg_op1[2]_9639 ), .B
       (\genblk2.pcpi_div_minus_2470_59_n_487 ), .Y (n_6533));
  OR2X1 g90318__5107(.A (mem_state[0]), .B (mem_state[1]), .Y (n_6050));
  NOR2BX1 g90319__6260(.AN (mem_wordsize[0]), .B (mem_wordsize[1]), .Y
       (n_5980));
  NOR2X1 g90321__4319(.A (instr_andi), .B (instr_and), .Y (n_6048));
  OR2X1 g90323__8428(.A (mem_wordsize[0]), .B (n_5993), .Y (n_5984));
  NOR2X2 g90324__5526(.A (mem_wordsize[0]), .B (mem_wordsize[1]), .Y
       (n_608));
  AND2X2 g90325__6783(.A (n_5995), .B (n_5994), .Y (n_5974));
  OR2X2 g90327__3680(.A (mem_do_prefetch), .B (mem_do_rinst), .Y
       (n_313));
  INVXL g90328(.A (mem_rdata[1]), .Y (n_6027));
  INVXL g90329(.A (latched_store), .Y (n_6026));
  INVX1 g90346(.A (mem_rdata[0]), .Y (n_6011));
  DFFX1 \genblk2.pcpi_div_pcpi_wait_reg (.CK (clk), .D (n_6290), .Q
       (pcpi_div_wait), .QN (n_5999));
  INVX2 drc_bufs90393(.A (n_120), .Y (n_119));
  INVX1 drc_bufs90399(.A (n_5984), .Y (n_5996));
  INVX3 drc_bufs90410(.A (n_320), .Y (n_5997));
  INVX1 drc_bufs90413(.A (n_608), .Y (n_6517));
  INVX1 drc_bufs90432(.A (n_5980), .Y (n_56));
  INVX1 drc_bufs90472(.A (n_48), .Y (n_5970));
  INVXL drc_bufs90481(.A (\genblk2.pcpi_div_n_2109 ), .Y (n_5995));
  INVX1 drc_bufs90513(.A (n_331), .Y (n_5998));
  INVX1 drc_bufs90645(.A (\reg_op2[5]_9674 ), .Y (n_756));
  INVX1 drc_bufs90681(.A (\reg_op2[3]_9672 ), .Y (n_725));
  INVX1 drc_bufs90821(.A (\reg_op1[4]_9641 ), .Y (n_717));
  INVX1 drc_bufs90825(.A (\reg_op1[5]_9642 ), .Y (n_5859));
  INVX1 drc_bufs90882(.A (\reg_op1[30]_9667 ), .Y (n_718));
  INVX1 drc_bufs90886(.A (\reg_op1[27]_9664 ), .Y (n_5829));
  INVX1 drc_bufs90890(.A (\reg_op1[23]_9660 ), .Y (n_5827));
  INVX1 drc_bufs90906(.A (\reg_op2[4]_9673 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_477 ));
  INVX1 drc_bufs90918(.A (\reg_op1[16]_9653 ), .Y (n_5813));
  INVX1 drc_bufs90922(.A (mem_wordsize[1]), .Y (n_5993));
  INVX1 drc_bufs90990(.A (\reg_op1[29]_9666 ), .Y (n_716));
  INVX1 drc_bufs90994(.A (\reg_op1[28]_9665 ), .Y (n_5788));
  INVX1 drc_bufs90998(.A (\reg_op1[26]_9663 ), .Y (n_5786));
  INVX1 drc_bufs91002(.A (\reg_op1[25]_9662 ), .Y (n_5784));
  INVX1 drc_bufs91006(.A (\reg_op1[24]_9661 ), .Y (n_713));
  INVX1 drc_bufs91010(.A (\reg_op1[17]_9654 ), .Y (n_715));
  INVX1 drc_bufs91014(.A (\reg_op1[20]_9657 ), .Y (n_634));
  OR2X1 g2__1617(.A (instr_or), .B (instr_ori), .Y (n_120));
  OR3X1 g91910__2802(.A (clear_prefetched_high_word_q), .B (n_6524), .C
       (n_6531), .Y (n_48));
  OR2X1 g91911__1705(.A (instr_xori), .B (instr_xor), .Y (n_279));
  NAND2X1 g91912__5122(.A (n_6060), .B (n_6287), .Y (mem_xfer));
  NOR2BX4 g91913__8246(.AN (n_5994), .B (n_5995), .Y (n_5694));
  DFFHQX1 \alu_out_q_reg[0] (.CK (clk), .D (n_5515), .Q (alu_out_q[0]));
  DFFHQX1 \alu_out_q_reg[1] (.CK (clk), .D (n_2281), .Q (alu_out_q[1]));
  DFFHQX1 \alu_out_q_reg[6] (.CK (clk), .D (n_2118), .Q (alu_out_q[6]));
  DFFHQX1 \alu_out_q_reg[7] (.CK (clk), .D (n_2119), .Q (alu_out_q[7]));
  DFFHQX1 \alu_out_q_reg[8] (.CK (clk), .D (n_2279), .Q (alu_out_q[8]));
  DFFHQX1 \alu_out_q_reg[9] (.CK (clk), .D (n_2280), .Q (alu_out_q[9]));
  DFFHQX1 \alu_out_q_reg[10] (.CK (clk), .D (n_2117), .Q
       (alu_out_q[10]));
  DFFHQX1 \alu_out_q_reg[11] (.CK (clk), .D (n_2121), .Q
       (alu_out_q[11]));
  DFFHQX1 \alu_out_q_reg[12] (.CK (clk), .D (n_2116), .Q
       (alu_out_q[12]));
  DFFHQX1 \alu_out_q_reg[13] (.CK (clk), .D (n_2122), .Q
       (alu_out_q[13]));
  DFFHQX1 \alu_out_q_reg[14] (.CK (clk), .D (n_2115), .Q
       (alu_out_q[14]));
  DFFHQX1 \alu_out_q_reg[15] (.CK (clk), .D (n_2120), .Q
       (alu_out_q[15]));
  DFFHQX1 \alu_out_q_reg[18] (.CK (clk), .D (n_2114), .Q
       (alu_out_q[18]));
  DFFHQX1 compressed_instr_reg(.CK (clk), .D (n_1555), .Q
       (compressed_instr));
  DFFHQX1 \count_cycle_reg[0] (.CK (clk), .D (n_896), .Q
       (count_cycle[0]));
  DFFHQX1 \count_cycle_reg[1] (.CK (clk), .D (n_800), .Q
       (count_cycle[1]));
  DFFHQX1 \count_cycle_reg[2] (.CK (clk), .D (n_946), .Q
       (count_cycle[2]));
  DFFHQX1 \count_cycle_reg[3] (.CK (clk), .D (n_794), .Q
       (count_cycle[3]));
  DFFHQX1 \count_cycle_reg[4] (.CK (clk), .D (n_925), .Q
       (count_cycle[4]));
  DFFHQX1 \count_cycle_reg[5] (.CK (clk), .D (n_948), .Q
       (count_cycle[5]));
  DFFHQX1 \count_cycle_reg[6] (.CK (clk), .D (n_799), .Q
       (count_cycle[6]));
  DFFHQX1 \count_cycle_reg[7] (.CK (clk), .D (n_796), .Q
       (count_cycle[7]));
  DFFHQX1 \count_cycle_reg[8] (.CK (clk), .D (n_813), .Q
       (count_cycle[8]));
  DFFHQX1 \count_cycle_reg[9] (.CK (clk), .D (n_795), .Q
       (count_cycle[9]));
  DFFHQX1 \count_cycle_reg[10] (.CK (clk), .D (n_950), .Q
       (count_cycle[10]));
  DFFHQX1 \count_cycle_reg[11] (.CK (clk), .D (n_894), .Q
       (count_cycle[11]));
  DFFHQX1 \count_cycle_reg[12] (.CK (clk), .D (n_924), .Q
       (count_cycle[12]));
  DFFHQX1 \count_cycle_reg[13] (.CK (clk), .D (n_939), .Q
       (count_cycle[13]));
  DFFHQX1 \count_cycle_reg[14] (.CK (clk), .D (n_898), .Q
       (count_cycle[14]));
  DFFHQX1 \count_cycle_reg[15] (.CK (clk), .D (n_888), .Q
       (count_cycle[15]));
  DFFHQX1 \count_cycle_reg[16] (.CK (clk), .D (n_818), .Q
       (count_cycle[16]));
  DFFHQX1 \count_cycle_reg[17] (.CK (clk), .D (n_951), .Q
       (count_cycle[17]));
  DFFHQX1 \count_cycle_reg[18] (.CK (clk), .D (n_826), .Q
       (count_cycle[18]));
  DFFHQX1 \count_cycle_reg[19] (.CK (clk), .D (n_910), .Q
       (count_cycle[19]));
  DFFHQX1 \count_cycle_reg[20] (.CK (clk), .D (n_902), .Q
       (count_cycle[20]));
  DFFHQX1 \count_cycle_reg[21] (.CK (clk), .D (n_808), .Q
       (count_cycle[21]));
  DFFHQX1 \count_cycle_reg[22] (.CK (clk), .D (n_943), .Q
       (count_cycle[22]));
  DFFHQX1 \count_cycle_reg[23] (.CK (clk), .D (n_822), .Q
       (count_cycle[23]));
  DFFHQX1 \count_cycle_reg[24] (.CK (clk), .D (n_938), .Q
       (count_cycle[24]));
  DFFHQX1 \count_cycle_reg[25] (.CK (clk), .D (n_927), .Q
       (count_cycle[25]));
  DFFHQX1 \count_cycle_reg[26] (.CK (clk), .D (n_918), .Q
       (count_cycle[26]));
  DFFHQX1 \count_cycle_reg[27] (.CK (clk), .D (n_782), .Q
       (count_cycle[27]));
  DFFHQX1 \count_cycle_reg[28] (.CK (clk), .D (n_889), .Q
       (count_cycle[28]));
  DFFHQX1 \count_cycle_reg[29] (.CK (clk), .D (n_895), .Q
       (count_cycle[29]));
  DFFHQX1 \count_cycle_reg[30] (.CK (clk), .D (n_806), .Q
       (count_cycle[30]));
  DFFHQX1 \count_cycle_reg[31] (.CK (clk), .D (n_893), .Q
       (count_cycle[31]));
  DFFHQX1 \count_cycle_reg[32] (.CK (clk), .D (n_899), .Q
       (count_cycle[32]));
  DFFHQX1 \count_cycle_reg[33] (.CK (clk), .D (n_802), .Q
       (count_cycle[33]));
  DFFHQX1 \count_cycle_reg[34] (.CK (clk), .D (n_922), .Q
       (count_cycle[34]));
  DFFHQX1 \count_cycle_reg[35] (.CK (clk), .D (n_933), .Q
       (count_cycle[35]));
  DFFHQX1 \count_cycle_reg[36] (.CK (clk), .D (n_904), .Q
       (count_cycle[36]));
  DFFHQX1 \count_cycle_reg[37] (.CK (clk), .D (n_817), .Q
       (count_cycle[37]));
  DFFHQX1 \count_cycle_reg[38] (.CK (clk), .D (n_920), .Q
       (count_cycle[38]));
  DFFHQX1 \count_cycle_reg[39] (.CK (clk), .D (n_919), .Q
       (count_cycle[39]));
  DFFHQX1 \count_cycle_reg[40] (.CK (clk), .D (n_908), .Q
       (count_cycle[40]));
  DFFHQX1 \count_cycle_reg[41] (.CK (clk), .D (n_934), .Q
       (count_cycle[41]));
  DFFHQX1 \count_cycle_reg[42] (.CK (clk), .D (n_797), .Q
       (count_cycle[42]));
  DFFHQX1 \count_cycle_reg[43] (.CK (clk), .D (n_830), .Q
       (count_cycle[43]));
  DFFHQX1 \count_cycle_reg[44] (.CK (clk), .D (n_783), .Q
       (count_cycle[44]));
  DFFHQX1 \count_cycle_reg[45] (.CK (clk), .D (n_944), .Q
       (count_cycle[45]));
  DFFHQX1 \count_cycle_reg[46] (.CK (clk), .D (n_815), .Q
       (count_cycle[46]));
  DFFHQX1 \count_cycle_reg[47] (.CK (clk), .D (n_932), .Q
       (count_cycle[47]));
  DFFHQX1 \count_cycle_reg[48] (.CK (clk), .D (n_801), .Q
       (count_cycle[48]));
  DFFHQX1 \count_cycle_reg[49] (.CK (clk), .D (n_886), .Q
       (count_cycle[49]));
  DFFHQX1 \count_cycle_reg[50] (.CK (clk), .D (n_912), .Q
       (count_cycle[50]));
  DFFHQX1 \count_cycle_reg[51] (.CK (clk), .D (n_909), .Q
       (count_cycle[51]));
  DFFHQX1 \count_cycle_reg[52] (.CK (clk), .D (n_913), .Q
       (count_cycle[52]));
  DFFHQX1 \count_cycle_reg[53] (.CK (clk), .D (n_784), .Q
       (count_cycle[53]));
  DFFHQX1 \count_cycle_reg[54] (.CK (clk), .D (n_929), .Q
       (count_cycle[54]));
  DFFHQX1 \count_cycle_reg[55] (.CK (clk), .D (n_941), .Q
       (count_cycle[55]));
  DFFHQX1 \count_cycle_reg[56] (.CK (clk), .D (n_814), .Q
       (count_cycle[56]));
  DFFHQX1 \count_cycle_reg[57] (.CK (clk), .D (n_829), .Q
       (count_cycle[57]));
  DFFHQX1 \count_cycle_reg[58] (.CK (clk), .D (n_790), .Q
       (count_cycle[58]));
  DFFHQX1 \count_cycle_reg[59] (.CK (clk), .D (n_811), .Q
       (count_cycle[59]));
  DFFHQX1 \count_cycle_reg[60] (.CK (clk), .D (n_926), .Q
       (count_cycle[60]));
  DFFHQX1 \count_cycle_reg[61] (.CK (clk), .D (n_928), .Q
       (count_cycle[61]));
  DFFHQX1 \count_cycle_reg[62] (.CK (clk), .D (n_891), .Q
       (count_cycle[62]));
  DFFHQX1 \count_cycle_reg[63] (.CK (clk), .D (n_907), .Q
       (count_cycle[63]));
  DFFHQX1 \count_instr_reg[0] (.CK (clk), .D (n_1917), .Q
       (count_instr[0]));
  DFFHQX1 \count_instr_reg[1] (.CK (clk), .D (n_1819), .Q
       (count_instr[1]));
  DFFHQX1 \count_instr_reg[2] (.CK (clk), .D (n_1864), .Q
       (count_instr[2]));
  DFFHQX1 \count_instr_reg[3] (.CK (clk), .D (n_1868), .Q
       (count_instr[3]));
  DFFHQX1 \count_instr_reg[4] (.CK (clk), .D (n_1902), .Q
       (count_instr[4]));
  DFFHQX1 \count_instr_reg[5] (.CK (clk), .D (n_1826), .Q
       (count_instr[5]));
  DFFHQX1 \count_instr_reg[6] (.CK (clk), .D (n_1870), .Q
       (count_instr[6]));
  DFFHQX1 \count_instr_reg[7] (.CK (clk), .D (n_1913), .Q
       (count_instr[7]));
  DFFHQX1 \count_instr_reg[8] (.CK (clk), .D (n_1829), .Q
       (count_instr[8]));
  DFFHQX1 \count_instr_reg[9] (.CK (clk), .D (n_1875), .Q
       (count_instr[9]));
  DFFHQX1 \count_instr_reg[10] (.CK (clk), .D (n_1885), .Q
       (count_instr[10]));
  DFFHQX1 \count_instr_reg[11] (.CK (clk), .D (n_1821), .Q
       (count_instr[11]));
  DFFHQX1 \count_instr_reg[12] (.CK (clk), .D (n_1909), .Q
       (count_instr[12]));
  DFFHQX1 \count_instr_reg[13] (.CK (clk), .D (n_1817), .Q
       (count_instr[13]));
  DFFHQX1 \count_instr_reg[14] (.CK (clk), .D (n_1820), .Q
       (count_instr[14]));
  DFFHQX1 \count_instr_reg[15] (.CK (clk), .D (n_1827), .Q
       (count_instr[15]));
  DFFHQX1 \count_instr_reg[16] (.CK (clk), .D (n_1861), .Q
       (count_instr[16]));
  DFFHQX1 \count_instr_reg[17] (.CK (clk), .D (n_1831), .Q
       (count_instr[17]));
  DFFHQX1 \count_instr_reg[18] (.CK (clk), .D (n_1905), .Q
       (count_instr[18]));
  DFFHQX1 \count_instr_reg[19] (.CK (clk), .D (n_1906), .Q
       (count_instr[19]));
  DFFHQX1 \count_instr_reg[20] (.CK (clk), .D (n_1904), .Q
       (count_instr[20]));
  DFFHQX1 \count_instr_reg[21] (.CK (clk), .D (n_1822), .Q
       (count_instr[21]));
  DFFHQX1 \count_instr_reg[22] (.CK (clk), .D (n_1907), .Q
       (count_instr[22]));
  DFFHQX1 \count_instr_reg[23] (.CK (clk), .D (n_1818), .Q
       (count_instr[23]));
  DFFHQX1 \count_instr_reg[24] (.CK (clk), .D (n_1908), .Q
       (count_instr[24]));
  DFFHQX1 \count_instr_reg[25] (.CK (clk), .D (n_1823), .Q
       (count_instr[25]));
  DFFHQX1 \count_instr_reg[26] (.CK (clk), .D (n_1911), .Q
       (count_instr[26]));
  DFFHQX1 \count_instr_reg[27] (.CK (clk), .D (n_1910), .Q
       (count_instr[27]));
  DFFHQX1 \count_instr_reg[28] (.CK (clk), .D (n_1824), .Q
       (count_instr[28]));
  DFFHQX1 \count_instr_reg[29] (.CK (clk), .D (n_1825), .Q
       (count_instr[29]));
  DFFHQX1 \count_instr_reg[30] (.CK (clk), .D (n_1830), .Q
       (count_instr[30]));
  DFFHQX1 \count_instr_reg[31] (.CK (clk), .D (n_1857), .Q
       (count_instr[31]));
  DFFHQX1 \count_instr_reg[32] (.CK (clk), .D (n_1860), .Q
       (count_instr[32]));
  DFFHQX1 \count_instr_reg[33] (.CK (clk), .D (n_1859), .Q
       (count_instr[33]));
  DFFHQX1 \count_instr_reg[34] (.CK (clk), .D (n_1912), .Q
       (count_instr[34]));
  DFFHQX1 \count_instr_reg[35] (.CK (clk), .D (n_1833), .Q
       (count_instr[35]));
  DFFHQX1 \count_instr_reg[36] (.CK (clk), .D (n_1858), .Q
       (count_instr[36]));
  DFFHQX1 \count_instr_reg[37] (.CK (clk), .D (n_1856), .Q
       (count_instr[37]));
  DFFHQX1 \count_instr_reg[38] (.CK (clk), .D (n_1865), .Q
       (count_instr[38]));
  DFFHQX1 \count_instr_reg[39] (.CK (clk), .D (n_1832), .Q
       (count_instr[39]));
  DFFHQX1 \count_instr_reg[40] (.CK (clk), .D (n_1872), .Q
       (count_instr[40]));
  DFFHQX1 \count_instr_reg[41] (.CK (clk), .D (n_1855), .Q
       (count_instr[41]));
  DFFHQX1 \count_instr_reg[42] (.CK (clk), .D (n_1854), .Q
       (count_instr[42]));
  DFFHQX1 \count_instr_reg[43] (.CK (clk), .D (n_1828), .Q
       (count_instr[43]));
  DFFHQX1 \count_instr_reg[44] (.CK (clk), .D (n_1852), .Q
       (count_instr[44]));
  DFFHQX1 \count_instr_reg[45] (.CK (clk), .D (n_1853), .Q
       (count_instr[45]));
  DFFHQX1 \count_instr_reg[46] (.CK (clk), .D (n_1851), .Q
       (count_instr[46]));
  DFFHQX1 \count_instr_reg[47] (.CK (clk), .D (n_1850), .Q
       (count_instr[47]));
  DFFHQX1 \count_instr_reg[48] (.CK (clk), .D (n_1849), .Q
       (count_instr[48]));
  DFFHQX1 \count_instr_reg[49] (.CK (clk), .D (n_1848), .Q
       (count_instr[49]));
  DFFHQX1 \count_instr_reg[50] (.CK (clk), .D (n_1845), .Q
       (count_instr[50]));
  DFFHQX1 \count_instr_reg[51] (.CK (clk), .D (n_1847), .Q
       (count_instr[51]));
  DFFHQX1 \count_instr_reg[52] (.CK (clk), .D (n_1846), .Q
       (count_instr[52]));
  DFFHQX1 \count_instr_reg[53] (.CK (clk), .D (n_1844), .Q
       (count_instr[53]));
  DFFHQX1 \count_instr_reg[54] (.CK (clk), .D (n_1843), .Q
       (count_instr[54]));
  DFFHQX1 \count_instr_reg[55] (.CK (clk), .D (n_1842), .Q
       (count_instr[55]));
  DFFHQX1 \count_instr_reg[56] (.CK (clk), .D (n_1841), .Q
       (count_instr[56]));
  DFFHQX1 \count_instr_reg[57] (.CK (clk), .D (n_1840), .Q
       (count_instr[57]));
  DFFHQX1 \count_instr_reg[58] (.CK (clk), .D (n_1839), .Q
       (count_instr[58]));
  DFFHQX1 \count_instr_reg[59] (.CK (clk), .D (n_1838), .Q
       (count_instr[59]));
  DFFHQX1 \count_instr_reg[60] (.CK (clk), .D (n_1837), .Q
       (count_instr[60]));
  DFFHQX1 \count_instr_reg[61] (.CK (clk), .D (n_1836), .Q
       (count_instr[61]));
  DFFHQX1 \count_instr_reg[62] (.CK (clk), .D (n_1835), .Q
       (count_instr[62]));
  DFFHQX1 \count_instr_reg[63] (.CK (clk), .D (n_1834), .Q
       (count_instr[63]));
  DFFHQX1 \cpu_state_reg[0] (.CK (clk), .D (n_5066), .Q (cpu_state[0]));
  DFFHQX1 \cpu_state_reg[1] (.CK (clk), .D (n_5064), .Q (cpu_state[1]));
  DFFHQX1 \cpu_state_reg[7] (.CK (clk), .D (n_5149), .Q (cpu_state[7]));
  DFFHQX1 \cpuregs_reg[1][0] (.CK (clk), .D (n_3135), .Q
       (\cpuregs[1] [0]));
  DFFHQX1 \cpuregs_reg[1][1] (.CK (clk), .D (n_3209), .Q
       (\cpuregs[1] [1]));
  DFFHQX1 \cpuregs_reg[1][2] (.CK (clk), .D (n_3210), .Q
       (\cpuregs[1] [2]));
  DFFHQX1 \cpuregs_reg[1][3] (.CK (clk), .D (n_3119), .Q
       (\cpuregs[1] [3]));
  DFFHQX1 \cpuregs_reg[1][4] (.CK (clk), .D (n_3164), .Q
       (\cpuregs[1] [4]));
  DFFHQX1 \cpuregs_reg[1][5] (.CK (clk), .D (n_3163), .Q
       (\cpuregs[1] [5]));
  DFFHQX1 \cpuregs_reg[1][6] (.CK (clk), .D (n_3162), .Q
       (\cpuregs[1] [6]));
  DFFHQX1 \cpuregs_reg[1][7] (.CK (clk), .D (n_3161), .Q
       (\cpuregs[1] [7]));
  DFFHQX1 \cpuregs_reg[1][8] (.CK (clk), .D (n_3160), .Q
       (\cpuregs[1] [8]));
  DFFHQX1 \cpuregs_reg[1][9] (.CK (clk), .D (n_3159), .Q
       (\cpuregs[1] [9]));
  DFFHQX1 \cpuregs_reg[1][10] (.CK (clk), .D (n_3158), .Q
       (\cpuregs[1] [10]));
  DFFHQX1 \cpuregs_reg[1][11] (.CK (clk), .D (n_3157), .Q
       (\cpuregs[1] [11]));
  DFFHQX1 \cpuregs_reg[1][12] (.CK (clk), .D (n_3153), .Q
       (\cpuregs[1] [12]));
  DFFHQX1 \cpuregs_reg[1][13] (.CK (clk), .D (n_3156), .Q
       (\cpuregs[1] [13]));
  DFFHQX1 \cpuregs_reg[1][14] (.CK (clk), .D (n_3155), .Q
       (\cpuregs[1] [14]));
  DFFHQX1 \cpuregs_reg[1][15] (.CK (clk), .D (n_3154), .Q
       (\cpuregs[1] [15]));
  DFFHQX1 \cpuregs_reg[1][16] (.CK (clk), .D (n_3152), .Q
       (\cpuregs[1] [16]));
  DFFHQX1 \cpuregs_reg[1][17] (.CK (clk), .D (n_3151), .Q
       (\cpuregs[1] [17]));
  DFFHQX1 \cpuregs_reg[1][18] (.CK (clk), .D (n_3150), .Q
       (\cpuregs[1] [18]));
  DFFHQX1 \cpuregs_reg[1][19] (.CK (clk), .D (n_3149), .Q
       (\cpuregs[1] [19]));
  DFFHQX1 \cpuregs_reg[1][20] (.CK (clk), .D (n_3148), .Q
       (\cpuregs[1] [20]));
  DFFHQX1 \cpuregs_reg[1][21] (.CK (clk), .D (n_3147), .Q
       (\cpuregs[1] [21]));
  DFFHQX1 \cpuregs_reg[1][22] (.CK (clk), .D (n_3146), .Q
       (\cpuregs[1] [22]));
  DFFHQX1 \cpuregs_reg[1][23] (.CK (clk), .D (n_3145), .Q
       (\cpuregs[1] [23]));
  DFFHQX1 \cpuregs_reg[1][24] (.CK (clk), .D (n_3143), .Q
       (\cpuregs[1] [24]));
  DFFHQX1 \cpuregs_reg[1][25] (.CK (clk), .D (n_3144), .Q
       (\cpuregs[1] [25]));
  DFFHQX1 \cpuregs_reg[1][26] (.CK (clk), .D (n_3142), .Q
       (\cpuregs[1] [26]));
  DFFHQX1 \cpuregs_reg[1][27] (.CK (clk), .D (n_3141), .Q
       (\cpuregs[1] [27]));
  DFFHQX1 \cpuregs_reg[1][28] (.CK (clk), .D (n_3140), .Q
       (\cpuregs[1] [28]));
  DFFHQX1 \cpuregs_reg[1][29] (.CK (clk), .D (n_3137), .Q
       (\cpuregs[1] [29]));
  DFFHQX1 \cpuregs_reg[1][30] (.CK (clk), .D (n_3139), .Q
       (\cpuregs[1] [30]));
  DFFHQX1 \cpuregs_reg[1][31] (.CK (clk), .D (n_3138), .Q
       (\cpuregs[1] [31]));
  DFFHQX1 \cpuregs_reg[2][0] (.CK (clk), .D (n_3571), .Q
       (\cpuregs[2] [0]));
  DFFHQX1 \cpuregs_reg[2][1] (.CK (clk), .D (n_3988), .Q
       (\cpuregs[2] [1]));
  DFFHQX1 \cpuregs_reg[2][2] (.CK (clk), .D (n_3985), .Q
       (\cpuregs[2] [2]));
  DFFHQX1 \cpuregs_reg[2][3] (.CK (clk), .D (n_3991), .Q
       (\cpuregs[2] [3]));
  DFFHQX1 \cpuregs_reg[2][4] (.CK (clk), .D (n_3982), .Q
       (\cpuregs[2] [4]));
  DFFHQX1 \cpuregs_reg[2][5] (.CK (clk), .D (n_3974), .Q
       (\cpuregs[2] [5]));
  DFFHQX1 \cpuregs_reg[2][6] (.CK (clk), .D (n_3980), .Q
       (\cpuregs[2] [6]));
  DFFHQX1 \cpuregs_reg[2][7] (.CK (clk), .D (n_3977), .Q
       (\cpuregs[2] [7]));
  DFFHQX1 \cpuregs_reg[2][8] (.CK (clk), .D (n_3972), .Q
       (\cpuregs[2] [8]));
  DFFHQX1 \cpuregs_reg[2][9] (.CK (clk), .D (n_3969), .Q
       (\cpuregs[2] [9]));
  DFFHQX1 \cpuregs_reg[2][10] (.CK (clk), .D (n_3966), .Q
       (\cpuregs[2] [10]));
  DFFHQX1 \cpuregs_reg[2][11] (.CK (clk), .D (n_3963), .Q
       (\cpuregs[2] [11]));
  DFFHQX1 \cpuregs_reg[2][12] (.CK (clk), .D (n_4102), .Q
       (\cpuregs[2] [12]));
  DFFHQX1 \cpuregs_reg[2][13] (.CK (clk), .D (n_4099), .Q
       (\cpuregs[2] [13]));
  DFFHQX1 \cpuregs_reg[2][14] (.CK (clk), .D (n_4103), .Q
       (\cpuregs[2] [14]));
  DFFHQX1 \cpuregs_reg[2][15] (.CK (clk), .D (n_4120), .Q
       (\cpuregs[2] [15]));
  DFFHQX1 \cpuregs_reg[2][16] (.CK (clk), .D (n_4124), .Q
       (\cpuregs[2] [16]));
  DFFHQX1 \cpuregs_reg[2][17] (.CK (clk), .D (n_4125), .Q
       (\cpuregs[2] [17]));
  DFFHQX1 \cpuregs_reg[2][18] (.CK (clk), .D (n_4130), .Q
       (\cpuregs[2] [18]));
  DFFHQX1 \cpuregs_reg[2][19] (.CK (clk), .D (n_4132), .Q
       (\cpuregs[2] [19]));
  DFFHQX1 \cpuregs_reg[2][20] (.CK (clk), .D (n_4134), .Q
       (\cpuregs[2] [20]));
  DFFHQX1 \cpuregs_reg[2][21] (.CK (clk), .D (n_4139), .Q
       (\cpuregs[2] [21]));
  DFFHQX1 \cpuregs_reg[2][22] (.CK (clk), .D (n_4140), .Q
       (\cpuregs[2] [22]));
  DFFHQX1 \cpuregs_reg[2][23] (.CK (clk), .D (n_4142), .Q
       (\cpuregs[2] [23]));
  DFFHQX1 \cpuregs_reg[2][24] (.CK (clk), .D (n_4153), .Q
       (\cpuregs[2] [24]));
  DFFHQX1 \cpuregs_reg[2][25] (.CK (clk), .D (n_4147), .Q
       (\cpuregs[2] [25]));
  DFFHQX1 \cpuregs_reg[2][26] (.CK (clk), .D (n_4151), .Q
       (\cpuregs[2] [26]));
  DFFHQX1 \cpuregs_reg[2][27] (.CK (clk), .D (n_4155), .Q
       (\cpuregs[2] [27]));
  DFFHQX1 \cpuregs_reg[2][28] (.CK (clk), .D (n_4157), .Q
       (\cpuregs[2] [28]));
  DFFHQX1 \cpuregs_reg[2][29] (.CK (clk), .D (n_4161), .Q
       (\cpuregs[2] [29]));
  DFFHQX1 \cpuregs_reg[2][30] (.CK (clk), .D (n_4164), .Q
       (\cpuregs[2] [30]));
  DFFHQX1 \cpuregs_reg[2][31] (.CK (clk), .D (n_4166), .Q
       (\cpuregs[2] [31]));
  DFFHQX1 \cpuregs_reg[3][0] (.CK (clk), .D (n_3569), .Q
       (\cpuregs[3] [0]));
  DFFHQX1 \cpuregs_reg[3][1] (.CK (clk), .D (n_4168), .Q
       (\cpuregs[3] [1]));
  DFFHQX1 \cpuregs_reg[3][2] (.CK (clk), .D (n_4169), .Q
       (\cpuregs[3] [2]));
  DFFHQX1 \cpuregs_reg[3][3] (.CK (clk), .D (n_4170), .Q
       (\cpuregs[3] [3]));
  DFFHQX1 \cpuregs_reg[3][4] (.CK (clk), .D (n_4175), .Q
       (\cpuregs[3] [4]));
  DFFHQX1 \cpuregs_reg[3][5] (.CK (clk), .D (n_4171), .Q
       (\cpuregs[3] [5]));
  DFFHQX1 \cpuregs_reg[3][6] (.CK (clk), .D (n_4172), .Q
       (\cpuregs[3] [6]));
  DFFHQX1 \cpuregs_reg[3][7] (.CK (clk), .D (n_4174), .Q
       (\cpuregs[3] [7]));
  DFFHQX1 \cpuregs_reg[3][8] (.CK (clk), .D (n_4176), .Q
       (\cpuregs[3] [8]));
  DFFHQX1 \cpuregs_reg[3][9] (.CK (clk), .D (n_4177), .Q
       (\cpuregs[3] [9]));
  DFFHQX1 \cpuregs_reg[3][10] (.CK (clk), .D (n_4178), .Q
       (\cpuregs[3] [10]));
  DFFHQX1 \cpuregs_reg[3][11] (.CK (clk), .D (n_4179), .Q
       (\cpuregs[3] [11]));
  DFFHQX1 \cpuregs_reg[3][12] (.CK (clk), .D (n_4180), .Q
       (\cpuregs[3] [12]));
  DFFHQX1 \cpuregs_reg[3][13] (.CK (clk), .D (n_4181), .Q
       (\cpuregs[3] [13]));
  DFFHQX1 \cpuregs_reg[3][14] (.CK (clk), .D (n_4183), .Q
       (\cpuregs[3] [14]));
  DFFHQX1 \cpuregs_reg[3][15] (.CK (clk), .D (n_4184), .Q
       (\cpuregs[3] [15]));
  DFFHQX1 \cpuregs_reg[3][16] (.CK (clk), .D (n_4188), .Q
       (\cpuregs[3] [16]));
  DFFHQX1 \cpuregs_reg[3][17] (.CK (clk), .D (n_4192), .Q
       (\cpuregs[3] [17]));
  DFFHQX1 \cpuregs_reg[3][18] (.CK (clk), .D (n_4194), .Q
       (\cpuregs[3] [18]));
  DFFHQX1 \cpuregs_reg[3][20] (.CK (clk), .D (n_4200), .Q
       (\cpuregs[3] [20]));
  DFFHQX1 \cpuregs_reg[3][23] (.CK (clk), .D (n_4209), .Q
       (\cpuregs[3] [23]));
  DFFHQX1 \cpuregs_reg[3][24] (.CK (clk), .D (n_4217), .Q
       (\cpuregs[3] [24]));
  DFFHQX1 \cpuregs_reg[3][25] (.CK (clk), .D (n_4214), .Q
       (\cpuregs[3] [25]));
  DFFHQX1 \cpuregs_reg[3][26] (.CK (clk), .D (n_4218), .Q
       (\cpuregs[3] [26]));
  DFFHQX1 \cpuregs_reg[3][27] (.CK (clk), .D (n_4222), .Q
       (\cpuregs[3] [27]));
  DFFHQX1 \cpuregs_reg[3][28] (.CK (clk), .D (n_4226), .Q
       (\cpuregs[3] [28]));
  DFFHQX1 \cpuregs_reg[3][29] (.CK (clk), .D (n_4227), .Q
       (\cpuregs[3] [29]));
  DFFHQX1 \cpuregs_reg[3][30] (.CK (clk), .D (n_4230), .Q
       (\cpuregs[3] [30]));
  DFFHQX1 \cpuregs_reg[3][31] (.CK (clk), .D (n_4232), .Q
       (\cpuregs[3] [31]));
  DFFHQX1 \cpuregs_reg[4][0] (.CK (clk), .D (n_3496), .Q
       (\cpuregs[4] [0]));
  DFFHQX1 \cpuregs_reg[4][1] (.CK (clk), .D (n_3760), .Q
       (\cpuregs[4] [1]));
  DFFHQX1 \cpuregs_reg[4][2] (.CK (clk), .D (n_3759), .Q
       (\cpuregs[4] [2]));
  DFFHQX1 \cpuregs_reg[4][3] (.CK (clk), .D (n_3758), .Q
       (\cpuregs[4] [3]));
  DFFHQX1 \cpuregs_reg[4][4] (.CK (clk), .D (n_3757), .Q
       (\cpuregs[4] [4]));
  DFFHQX1 \cpuregs_reg[4][5] (.CK (clk), .D (n_3755), .Q
       (\cpuregs[4] [5]));
  DFFHQX1 \cpuregs_reg[4][6] (.CK (clk), .D (n_3756), .Q
       (\cpuregs[4] [6]));
  DFFHQX1 \cpuregs_reg[4][7] (.CK (clk), .D (n_3754), .Q
       (\cpuregs[4] [7]));
  DFFHQX1 \cpuregs_reg[4][8] (.CK (clk), .D (n_3753), .Q
       (\cpuregs[4] [8]));
  DFFHQX1 \cpuregs_reg[4][9] (.CK (clk), .D (n_3752), .Q
       (\cpuregs[4] [9]));
  DFFHQX1 \cpuregs_reg[4][10] (.CK (clk), .D (n_3751), .Q
       (\cpuregs[4] [10]));
  DFFHQX1 \cpuregs_reg[4][11] (.CK (clk), .D (n_3750), .Q
       (\cpuregs[4] [11]));
  DFFHQX1 \cpuregs_reg[4][12] (.CK (clk), .D (n_3749), .Q
       (\cpuregs[4] [12]));
  DFFHQX1 \cpuregs_reg[4][13] (.CK (clk), .D (n_3748), .Q
       (\cpuregs[4] [13]));
  DFFHQX1 \cpuregs_reg[4][14] (.CK (clk), .D (n_3747), .Q
       (\cpuregs[4] [14]));
  DFFHQX1 \cpuregs_reg[4][15] (.CK (clk), .D (n_3746), .Q
       (\cpuregs[4] [15]));
  DFFHQX1 \cpuregs_reg[4][16] (.CK (clk), .D (n_3745), .Q
       (\cpuregs[4] [16]));
  DFFHQX1 \cpuregs_reg[4][17] (.CK (clk), .D (n_3743), .Q
       (\cpuregs[4] [17]));
  DFFHQX1 \cpuregs_reg[4][18] (.CK (clk), .D (n_3744), .Q
       (\cpuregs[4] [18]));
  DFFHQX1 \cpuregs_reg[4][19] (.CK (clk), .D (n_3742), .Q
       (\cpuregs[4] [19]));
  DFFHQX1 \cpuregs_reg[4][20] (.CK (clk), .D (n_3741), .Q
       (\cpuregs[4] [20]));
  DFFHQX1 \cpuregs_reg[4][21] (.CK (clk), .D (n_3740), .Q
       (\cpuregs[4] [21]));
  DFFHQX1 \cpuregs_reg[4][22] (.CK (clk), .D (n_3739), .Q
       (\cpuregs[4] [22]));
  DFFHQX1 \cpuregs_reg[4][23] (.CK (clk), .D (n_3738), .Q
       (\cpuregs[4] [23]));
  DFFHQX1 \cpuregs_reg[4][24] (.CK (clk), .D (n_3737), .Q
       (\cpuregs[4] [24]));
  DFFHQX1 \cpuregs_reg[4][25] (.CK (clk), .D (n_3736), .Q
       (\cpuregs[4] [25]));
  DFFHQX1 \cpuregs_reg[4][26] (.CK (clk), .D (n_3735), .Q
       (\cpuregs[4] [26]));
  DFFHQX1 \cpuregs_reg[4][27] (.CK (clk), .D (n_3734), .Q
       (\cpuregs[4] [27]));
  DFFHQX1 \cpuregs_reg[4][28] (.CK (clk), .D (n_3733), .Q
       (\cpuregs[4] [28]));
  DFFHQX1 \cpuregs_reg[4][29] (.CK (clk), .D (n_3732), .Q
       (\cpuregs[4] [29]));
  DFFHQX1 \cpuregs_reg[4][30] (.CK (clk), .D (n_3731), .Q
       (\cpuregs[4] [30]));
  DFFHQX1 \cpuregs_reg[4][31] (.CK (clk), .D (n_3730), .Q
       (\cpuregs[4] [31]));
  DFFHQX1 \cpuregs_reg[5][0] (.CK (clk), .D (n_3566), .Q
       (\cpuregs[5] [0]));
  DFFHQX1 \cpuregs_reg[5][1] (.CK (clk), .D (n_4266), .Q
       (\cpuregs[5] [1]));
  DFFHQX1 \cpuregs_reg[5][2] (.CK (clk), .D (n_4267), .Q
       (\cpuregs[5] [2]));
  DFFHQX1 \cpuregs_reg[5][3] (.CK (clk), .D (n_4268), .Q
       (\cpuregs[5] [3]));
  DFFHQX1 \cpuregs_reg[5][4] (.CK (clk), .D (n_4269), .Q
       (\cpuregs[5] [4]));
  DFFHQX1 \cpuregs_reg[5][5] (.CK (clk), .D (n_4270), .Q
       (\cpuregs[5] [5]));
  DFFHQX1 \cpuregs_reg[5][6] (.CK (clk), .D (n_4271), .Q
       (\cpuregs[5] [6]));
  DFFHQX1 \cpuregs_reg[5][7] (.CK (clk), .D (n_4272), .Q
       (\cpuregs[5] [7]));
  DFFHQX1 \cpuregs_reg[5][8] (.CK (clk), .D (n_4273), .Q
       (\cpuregs[5] [8]));
  DFFHQX1 \cpuregs_reg[5][9] (.CK (clk), .D (n_4274), .Q
       (\cpuregs[5] [9]));
  DFFHQX1 \cpuregs_reg[5][10] (.CK (clk), .D (n_4275), .Q
       (\cpuregs[5] [10]));
  DFFHQX1 \cpuregs_reg[5][11] (.CK (clk), .D (n_4276), .Q
       (\cpuregs[5] [11]));
  DFFHQX1 \cpuregs_reg[5][12] (.CK (clk), .D (n_4277), .Q
       (\cpuregs[5] [12]));
  DFFHQX1 \cpuregs_reg[5][13] (.CK (clk), .D (n_4278), .Q
       (\cpuregs[5] [13]));
  DFFHQX1 \cpuregs_reg[5][14] (.CK (clk), .D (n_4279), .Q
       (\cpuregs[5] [14]));
  DFFHQX1 \cpuregs_reg[5][15] (.CK (clk), .D (n_4280), .Q
       (\cpuregs[5] [15]));
  DFFHQX1 \cpuregs_reg[5][16] (.CK (clk), .D (n_4281), .Q
       (\cpuregs[5] [16]));
  DFFHQX1 \cpuregs_reg[5][17] (.CK (clk), .D (n_3715), .Q
       (\cpuregs[5] [17]));
  DFFHQX1 \cpuregs_reg[5][18] (.CK (clk), .D (n_3961), .Q
       (\cpuregs[5] [18]));
  DFFHQX1 \cpuregs_reg[5][19] (.CK (clk), .D (n_3960), .Q
       (\cpuregs[5] [19]));
  DFFHQX1 \cpuregs_reg[5][20] (.CK (clk), .D (n_3959), .Q
       (\cpuregs[5] [20]));
  DFFHQX1 \cpuregs_reg[5][21] (.CK (clk), .D (n_3958), .Q
       (\cpuregs[5] [21]));
  DFFHQX1 \cpuregs_reg[5][22] (.CK (clk), .D (n_3956), .Q
       (\cpuregs[5] [22]));
  DFFHQX1 \cpuregs_reg[5][23] (.CK (clk), .D (n_3957), .Q
       (\cpuregs[5] [23]));
  DFFHQX1 \cpuregs_reg[5][24] (.CK (clk), .D (n_3954), .Q
       (\cpuregs[5] [24]));
  DFFHQX1 \cpuregs_reg[5][25] (.CK (clk), .D (n_3953), .Q
       (\cpuregs[5] [25]));
  DFFHQX1 \cpuregs_reg[5][26] (.CK (clk), .D (n_3952), .Q
       (\cpuregs[5] [26]));
  DFFHQX1 \cpuregs_reg[5][27] (.CK (clk), .D (n_3951), .Q
       (\cpuregs[5] [27]));
  DFFHQX1 \cpuregs_reg[5][28] (.CK (clk), .D (n_3950), .Q
       (\cpuregs[5] [28]));
  DFFHQX1 \cpuregs_reg[5][29] (.CK (clk), .D (n_3949), .Q
       (\cpuregs[5] [29]));
  DFFHQX1 \cpuregs_reg[5][30] (.CK (clk), .D (n_3948), .Q
       (\cpuregs[5] [30]));
  DFFHQX1 \cpuregs_reg[5][31] (.CK (clk), .D (n_3946), .Q
       (\cpuregs[5] [31]));
  DFFHQX1 \cpuregs_reg[6][0] (.CK (clk), .D (n_3564), .Q
       (\cpuregs[6] [0]));
  DFFHQX1 \cpuregs_reg[6][1] (.CK (clk), .D (n_4265), .Q
       (\cpuregs[6] [1]));
  DFFHQX1 \cpuregs_reg[6][2] (.CK (clk), .D (n_4264), .Q
       (\cpuregs[6] [2]));
  DFFHQX1 \cpuregs_reg[6][3] (.CK (clk), .D (n_3936), .Q
       (\cpuregs[6] [3]));
  DFFHQX1 \cpuregs_reg[6][4] (.CK (clk), .D (n_3931), .Q
       (\cpuregs[6] [4]));
  DFFHQX1 \cpuregs_reg[6][5] (.CK (clk), .D (n_3930), .Q
       (\cpuregs[6] [5]));
  DFFHQX1 \cpuregs_reg[6][6] (.CK (clk), .D (n_3926), .Q
       (\cpuregs[6] [6]));
  DFFHQX1 \cpuregs_reg[6][7] (.CK (clk), .D (n_3924), .Q
       (\cpuregs[6] [7]));
  DFFHQX1 \cpuregs_reg[6][8] (.CK (clk), .D (n_3920), .Q
       (\cpuregs[6] [8]));
  DFFHQX1 \cpuregs_reg[6][9] (.CK (clk), .D (n_3917), .Q
       (\cpuregs[6] [9]));
  DFFHQX1 \cpuregs_reg[6][10] (.CK (clk), .D (n_3915), .Q
       (\cpuregs[6] [10]));
  DFFHQX1 \cpuregs_reg[6][11] (.CK (clk), .D (n_3913), .Q
       (\cpuregs[6] [11]));
  DFFHQX1 \cpuregs_reg[6][12] (.CK (clk), .D (n_3909), .Q
       (\cpuregs[6] [12]));
  DFFHQX1 \cpuregs_reg[6][13] (.CK (clk), .D (n_3906), .Q
       (\cpuregs[6] [13]));
  DFFHQX1 \cpuregs_reg[6][14] (.CK (clk), .D (n_3904), .Q
       (\cpuregs[6] [14]));
  DFFHQX1 \cpuregs_reg[6][15] (.CK (clk), .D (n_3902), .Q
       (\cpuregs[6] [15]));
  DFFHQX1 \cpuregs_reg[6][16] (.CK (clk), .D (n_3893), .Q
       (\cpuregs[6] [16]));
  DFFHQX1 \cpuregs_reg[6][17] (.CK (clk), .D (n_3899), .Q
       (\cpuregs[6] [17]));
  DFFHQX1 \cpuregs_reg[6][18] (.CK (clk), .D (n_3896), .Q
       (\cpuregs[6] [18]));
  DFFHQX1 \cpuregs_reg[6][19] (.CK (clk), .D (n_3891), .Q
       (\cpuregs[6] [19]));
  DFFHQX1 \cpuregs_reg[6][20] (.CK (clk), .D (n_3887), .Q
       (\cpuregs[6] [20]));
  DFFHQX1 \cpuregs_reg[6][21] (.CK (clk), .D (n_3886), .Q
       (\cpuregs[6] [21]));
  DFFHQX1 \cpuregs_reg[6][22] (.CK (clk), .D (n_3885), .Q
       (\cpuregs[6] [22]));
  DFFHQX1 \cpuregs_reg[6][23] (.CK (clk), .D (n_3883), .Q
       (\cpuregs[6] [23]));
  DFFHQX1 \cpuregs_reg[6][24] (.CK (clk), .D (n_3879), .Q
       (\cpuregs[6] [24]));
  DFFHQX1 \cpuregs_reg[6][25] (.CK (clk), .D (n_3874), .Q
       (\cpuregs[6] [25]));
  DFFHQX1 \cpuregs_reg[6][26] (.CK (clk), .D (n_3998), .Q
       (\cpuregs[6] [26]));
  DFFHQX1 \cpuregs_reg[6][27] (.CK (clk), .D (n_3872), .Q
       (\cpuregs[6] [27]));
  DFFHQX1 \cpuregs_reg[6][28] (.CK (clk), .D (n_3865), .Q
       (\cpuregs[6] [28]));
  DFFHQX1 \cpuregs_reg[6][29] (.CK (clk), .D (n_3863), .Q
       (\cpuregs[6] [29]));
  DFFHQX1 \cpuregs_reg[6][30] (.CK (clk), .D (n_3864), .Q
       (\cpuregs[6] [30]));
  DFFHQX1 \cpuregs_reg[6][31] (.CK (clk), .D (n_3862), .Q
       (\cpuregs[6] [31]));
  DFFHQX1 \cpuregs_reg[7][0] (.CK (clk), .D (n_3494), .Q
       (\cpuregs[7] [0]));
  DFFHQX1 \cpuregs_reg[7][1] (.CK (clk), .D (n_3729), .Q
       (\cpuregs[7] [1]));
  DFFHQX1 \cpuregs_reg[7][2] (.CK (clk), .D (n_3726), .Q
       (\cpuregs[7] [2]));
  DFFHQX1 \cpuregs_reg[7][3] (.CK (clk), .D (n_3728), .Q
       (\cpuregs[7] [3]));
  DFFHQX1 \cpuregs_reg[7][4] (.CK (clk), .D (n_3727), .Q
       (\cpuregs[7] [4]));
  DFFHQX1 \cpuregs_reg[7][5] (.CK (clk), .D (n_3725), .Q
       (\cpuregs[7] [5]));
  DFFHQX1 \cpuregs_reg[7][6] (.CK (clk), .D (n_3724), .Q
       (\cpuregs[7] [6]));
  DFFHQX1 \cpuregs_reg[7][7] (.CK (clk), .D (n_3723), .Q
       (\cpuregs[7] [7]));
  DFFHQX1 \cpuregs_reg[7][8] (.CK (clk), .D (n_3722), .Q
       (\cpuregs[7] [8]));
  DFFHQX1 \cpuregs_reg[7][9] (.CK (clk), .D (n_3721), .Q
       (\cpuregs[7] [9]));
  DFFHQX1 \cpuregs_reg[7][10] (.CK (clk), .D (n_3720), .Q
       (\cpuregs[7] [10]));
  DFFHQX1 \cpuregs_reg[7][11] (.CK (clk), .D (n_3719), .Q
       (\cpuregs[7] [11]));
  DFFHQX1 \cpuregs_reg[7][12] (.CK (clk), .D (n_3718), .Q
       (\cpuregs[7] [12]));
  DFFHQX1 \cpuregs_reg[7][13] (.CK (clk), .D (n_3717), .Q
       (\cpuregs[7] [13]));
  DFFHQX1 \cpuregs_reg[7][14] (.CK (clk), .D (n_3716), .Q
       (\cpuregs[7] [14]));
  DFFHQX1 \cpuregs_reg[7][15] (.CK (clk), .D (n_3962), .Q
       (\cpuregs[7] [15]));
  DFFHQX1 \cpuregs_reg[7][16] (.CK (clk), .D (n_3714), .Q
       (\cpuregs[7] [16]));
  DFFHQX1 \cpuregs_reg[7][17] (.CK (clk), .D (n_3713), .Q
       (\cpuregs[7] [17]));
  DFFHQX1 \cpuregs_reg[7][18] (.CK (clk), .D (n_3712), .Q
       (\cpuregs[7] [18]));
  DFFHQX1 \cpuregs_reg[7][19] (.CK (clk), .D (n_3711), .Q
       (\cpuregs[7] [19]));
  DFFHQX1 \cpuregs_reg[7][20] (.CK (clk), .D (n_3710), .Q
       (\cpuregs[7] [20]));
  DFFHQX1 \cpuregs_reg[7][21] (.CK (clk), .D (n_3709), .Q
       (\cpuregs[7] [21]));
  DFFHQX1 \cpuregs_reg[7][22] (.CK (clk), .D (n_3708), .Q
       (\cpuregs[7] [22]));
  DFFHQX1 \cpuregs_reg[7][23] (.CK (clk), .D (n_3707), .Q
       (\cpuregs[7] [23]));
  DFFHQX1 \cpuregs_reg[7][24] (.CK (clk), .D (n_3706), .Q
       (\cpuregs[7] [24]));
  DFFHQX1 \cpuregs_reg[7][25] (.CK (clk), .D (n_3705), .Q
       (\cpuregs[7] [25]));
  DFFHQX1 \cpuregs_reg[7][26] (.CK (clk), .D (n_3704), .Q
       (\cpuregs[7] [26]));
  DFFHQX1 \cpuregs_reg[7][27] (.CK (clk), .D (n_3703), .Q
       (\cpuregs[7] [27]));
  DFFHQX1 \cpuregs_reg[7][28] (.CK (clk), .D (n_3702), .Q
       (\cpuregs[7] [28]));
  DFFHQX1 \cpuregs_reg[7][29] (.CK (clk), .D (n_3701), .Q
       (\cpuregs[7] [29]));
  DFFHQX1 \cpuregs_reg[7][30] (.CK (clk), .D (n_3700), .Q
       (\cpuregs[7] [30]));
  DFFHQX1 \cpuregs_reg[7][31] (.CK (clk), .D (n_3699), .Q
       (\cpuregs[7] [31]));
  DFFHQX1 \cpuregs_reg[8][0] (.CK (clk), .D (n_3136), .Q
       (\cpuregs[8] [0]));
  DFFHQX1 \cpuregs_reg[8][1] (.CK (clk), .D (n_3178), .Q
       (\cpuregs[8] [1]));
  DFFHQX1 \cpuregs_reg[8][2] (.CK (clk), .D (n_3184), .Q
       (\cpuregs[8] [2]));
  DFFHQX1 \cpuregs_reg[8][3] (.CK (clk), .D (n_3179), .Q
       (\cpuregs[8] [3]));
  DFFHQX1 \cpuregs_reg[8][4] (.CK (clk), .D (n_3180), .Q
       (\cpuregs[8] [4]));
  DFFHQX1 \cpuregs_reg[8][5] (.CK (clk), .D (n_3181), .Q
       (\cpuregs[8] [5]));
  DFFHQX1 \cpuregs_reg[8][6] (.CK (clk), .D (n_3182), .Q
       (\cpuregs[8] [6]));
  DFFHQX1 \cpuregs_reg[8][7] (.CK (clk), .D (n_3183), .Q
       (\cpuregs[8] [7]));
  DFFHQX1 \cpuregs_reg[8][8] (.CK (clk), .D (n_3177), .Q
       (\cpuregs[8] [8]));
  DFFHQX1 \cpuregs_reg[8][9] (.CK (clk), .D (n_3186), .Q
       (\cpuregs[8] [9]));
  DFFHQX1 \cpuregs_reg[8][10] (.CK (clk), .D (n_3185), .Q
       (\cpuregs[8] [10]));
  DFFHQX1 \cpuregs_reg[8][11] (.CK (clk), .D (n_3187), .Q
       (\cpuregs[8] [11]));
  DFFHQX1 \cpuregs_reg[8][12] (.CK (clk), .D (n_3188), .Q
       (\cpuregs[8] [12]));
  DFFHQX1 \cpuregs_reg[8][13] (.CK (clk), .D (n_3189), .Q
       (\cpuregs[8] [13]));
  DFFHQX1 \cpuregs_reg[8][14] (.CK (clk), .D (n_3190), .Q
       (\cpuregs[8] [14]));
  DFFHQX1 \cpuregs_reg[8][15] (.CK (clk), .D (n_3192), .Q
       (\cpuregs[8] [15]));
  DFFHQX1 \cpuregs_reg[8][16] (.CK (clk), .D (n_3191), .Q
       (\cpuregs[8] [16]));
  DFFHQX1 \cpuregs_reg[8][17] (.CK (clk), .D (n_3194), .Q
       (\cpuregs[8] [17]));
  DFFHQX1 \cpuregs_reg[8][18] (.CK (clk), .D (n_3195), .Q
       (\cpuregs[8] [18]));
  DFFHQX1 \cpuregs_reg[8][19] (.CK (clk), .D (n_3196), .Q
       (\cpuregs[8] [19]));
  DFFHQX1 \cpuregs_reg[8][20] (.CK (clk), .D (n_3197), .Q
       (\cpuregs[8] [20]));
  DFFHQX1 \cpuregs_reg[8][21] (.CK (clk), .D (n_3200), .Q
       (\cpuregs[8] [21]));
  DFFHQX1 \cpuregs_reg[8][22] (.CK (clk), .D (n_3198), .Q
       (\cpuregs[8] [22]));
  DFFHQX1 \cpuregs_reg[8][23] (.CK (clk), .D (n_3199), .Q
       (\cpuregs[8] [23]));
  DFFHQX1 \cpuregs_reg[8][24] (.CK (clk), .D (n_3201), .Q
       (\cpuregs[8] [24]));
  DFFHQX1 \cpuregs_reg[8][25] (.CK (clk), .D (n_3202), .Q
       (\cpuregs[8] [25]));
  DFFHQX1 \cpuregs_reg[8][26] (.CK (clk), .D (n_3203), .Q
       (\cpuregs[8] [26]));
  DFFHQX1 \cpuregs_reg[8][27] (.CK (clk), .D (n_3204), .Q
       (\cpuregs[8] [27]));
  DFFHQX1 \cpuregs_reg[8][28] (.CK (clk), .D (n_3205), .Q
       (\cpuregs[8] [28]));
  DFFHQX1 \cpuregs_reg[8][29] (.CK (clk), .D (n_3206), .Q
       (\cpuregs[8] [29]));
  DFFHQX1 \cpuregs_reg[8][30] (.CK (clk), .D (n_3207), .Q
       (\cpuregs[8] [30]));
  DFFHQX1 \cpuregs_reg[8][31] (.CK (clk), .D (n_3208), .Q
       (\cpuregs[8] [31]));
  DFFHQX1 \cpuregs_reg[9][0] (.CK (clk), .D (n_3327), .Q
       (\cpuregs[9] [0]));
  DFFHQX1 \cpuregs_reg[9][1] (.CK (clk), .D (n_3409), .Q
       (\cpuregs[9] [1]));
  DFFHQX1 \cpuregs_reg[9][2] (.CK (clk), .D (n_3408), .Q
       (\cpuregs[9] [2]));
  DFFHQX1 \cpuregs_reg[9][3] (.CK (clk), .D (n_3406), .Q
       (\cpuregs[9] [3]));
  DFFHQX1 \cpuregs_reg[9][4] (.CK (clk), .D (n_3407), .Q
       (\cpuregs[9] [4]));
  DFFHQX1 \cpuregs_reg[9][5] (.CK (clk), .D (n_3405), .Q
       (\cpuregs[9] [5]));
  DFFHQX1 \cpuregs_reg[9][6] (.CK (clk), .D (n_3404), .Q
       (\cpuregs[9] [6]));
  DFFHQX1 \cpuregs_reg[9][7] (.CK (clk), .D (n_3403), .Q
       (\cpuregs[9] [7]));
  DFFHQX1 \cpuregs_reg[9][8] (.CK (clk), .D (n_3400), .Q
       (\cpuregs[9] [8]));
  DFFHQX1 \cpuregs_reg[9][9] (.CK (clk), .D (n_3402), .Q
       (\cpuregs[9] [9]));
  DFFHQX1 \cpuregs_reg[9][10] (.CK (clk), .D (n_3401), .Q
       (\cpuregs[9] [10]));
  DFFHQX1 \cpuregs_reg[9][11] (.CK (clk), .D (n_3399), .Q
       (\cpuregs[9] [11]));
  DFFHQX1 \cpuregs_reg[9][12] (.CK (clk), .D (n_3398), .Q
       (\cpuregs[9] [12]));
  DFFHQX1 \cpuregs_reg[9][13] (.CK (clk), .D (n_3397), .Q
       (\cpuregs[9] [13]));
  DFFHQX1 \cpuregs_reg[9][14] (.CK (clk), .D (n_3410), .Q
       (\cpuregs[9] [14]));
  DFFHQX1 \cpuregs_reg[9][15] (.CK (clk), .D (n_3417), .Q
       (\cpuregs[9] [15]));
  DFFHQX1 \cpuregs_reg[9][16] (.CK (clk), .D (n_3416), .Q
       (\cpuregs[9] [16]));
  DFFHQX1 \cpuregs_reg[9][17] (.CK (clk), .D (n_3423), .Q
       (\cpuregs[9] [17]));
  DFFHQX1 \cpuregs_reg[9][18] (.CK (clk), .D (n_3420), .Q
       (\cpuregs[9] [18]));
  DFFHQX1 \cpuregs_reg[9][19] (.CK (clk), .D (n_3421), .Q
       (\cpuregs[9] [19]));
  DFFHQX1 \cpuregs_reg[9][20] (.CK (clk), .D (n_3422), .Q
       (\cpuregs[9] [20]));
  DFFHQX1 \cpuregs_reg[9][21] (.CK (clk), .D (n_3428), .Q
       (\cpuregs[9] [21]));
  DFFHQX1 \cpuregs_reg[9][22] (.CK (clk), .D (n_3426), .Q
       (\cpuregs[9] [22]));
  DFFHQX1 \cpuregs_reg[9][23] (.CK (clk), .D (n_3427), .Q
       (\cpuregs[9] [23]));
  DFFHQX1 \cpuregs_reg[9][24] (.CK (clk), .D (n_3431), .Q
       (\cpuregs[9] [24]));
  DFFHQX1 \cpuregs_reg[9][25] (.CK (clk), .D (n_3432), .Q
       (\cpuregs[9] [25]));
  DFFHQX1 \cpuregs_reg[9][26] (.CK (clk), .D (n_3433), .Q
       (\cpuregs[9] [26]));
  DFFHQX1 \cpuregs_reg[9][27] (.CK (clk), .D (n_3393), .Q
       (\cpuregs[9] [27]));
  DFFHQX1 \cpuregs_reg[9][28] (.CK (clk), .D (n_3254), .Q
       (\cpuregs[9] [28]));
  DFFHQX1 \cpuregs_reg[9][29] (.CK (clk), .D (n_3394), .Q
       (\cpuregs[9] [29]));
  DFFHQX1 \cpuregs_reg[9][30] (.CK (clk), .D (n_3392), .Q
       (\cpuregs[9] [30]));
  DFFHQX1 \cpuregs_reg[9][31] (.CK (clk), .D (n_3391), .Q
       (\cpuregs[9] [31]));
  DFFHQX1 \cpuregs_reg[10][0] (.CK (clk), .D (n_3562), .Q
       (\cpuregs[10] [0]));
  DFFHQX1 \cpuregs_reg[10][1] (.CK (clk), .D (n_3859), .Q
       (\cpuregs[10] [1]));
  DFFHQX1 \cpuregs_reg[10][2] (.CK (clk), .D (n_3858), .Q
       (\cpuregs[10] [2]));
  DFFHQX1 \cpuregs_reg[10][3] (.CK (clk), .D (n_3860), .Q
       (\cpuregs[10] [3]));
  DFFHQX1 \cpuregs_reg[10][4] (.CK (clk), .D (n_3857), .Q
       (\cpuregs[10] [4]));
  DFFHQX1 \cpuregs_reg[10][5] (.CK (clk), .D (n_3856), .Q
       (\cpuregs[10] [5]));
  DFFHQX1 \cpuregs_reg[10][6] (.CK (clk), .D (n_3855), .Q
       (\cpuregs[10] [6]));
  DFFHQX1 \cpuregs_reg[10][7] (.CK (clk), .D (n_3854), .Q
       (\cpuregs[10] [7]));
  DFFHQX1 \cpuregs_reg[10][8] (.CK (clk), .D (n_3853), .Q
       (\cpuregs[10] [8]));
  DFFHQX1 \cpuregs_reg[10][9] (.CK (clk), .D (n_3852), .Q
       (\cpuregs[10] [9]));
  DFFHQX1 \cpuregs_reg[10][10] (.CK (clk), .D (n_3851), .Q
       (\cpuregs[10] [10]));
  DFFHQX1 \cpuregs_reg[10][11] (.CK (clk), .D (n_3850), .Q
       (\cpuregs[10] [11]));
  DFFHQX1 \cpuregs_reg[10][12] (.CK (clk), .D (n_3849), .Q
       (\cpuregs[10] [12]));
  DFFHQX1 \cpuregs_reg[10][13] (.CK (clk), .D (n_3848), .Q
       (\cpuregs[10] [13]));
  DFFHQX1 \cpuregs_reg[10][14] (.CK (clk), .D (n_3847), .Q
       (\cpuregs[10] [14]));
  DFFHQX1 \cpuregs_reg[10][15] (.CK (clk), .D (n_3845), .Q
       (\cpuregs[10] [15]));
  DFFHQX1 \cpuregs_reg[10][16] (.CK (clk), .D (n_3846), .Q
       (\cpuregs[10] [16]));
  DFFHQX1 \cpuregs_reg[10][17] (.CK (clk), .D (n_3844), .Q
       (\cpuregs[10] [17]));
  DFFHQX1 \cpuregs_reg[10][18] (.CK (clk), .D (n_3843), .Q
       (\cpuregs[10] [18]));
  DFFHQX1 \cpuregs_reg[10][19] (.CK (clk), .D (n_3842), .Q
       (\cpuregs[10] [19]));
  DFFHQX1 \cpuregs_reg[10][20] (.CK (clk), .D (n_3841), .Q
       (\cpuregs[10] [20]));
  DFFHQX1 \cpuregs_reg[10][21] (.CK (clk), .D (n_3839), .Q
       (\cpuregs[10] [21]));
  DFFHQX1 \cpuregs_reg[10][22] (.CK (clk), .D (n_3840), .Q
       (\cpuregs[10] [22]));
  DFFHQX1 \cpuregs_reg[10][23] (.CK (clk), .D (n_3838), .Q
       (\cpuregs[10] [23]));
  DFFHQX1 \cpuregs_reg[10][24] (.CK (clk), .D (n_3837), .Q
       (\cpuregs[10] [24]));
  DFFHQX1 \cpuregs_reg[10][25] (.CK (clk), .D (n_3836), .Q
       (\cpuregs[10] [25]));
  DFFHQX1 \cpuregs_reg[10][26] (.CK (clk), .D (n_3835), .Q
       (\cpuregs[10] [26]));
  DFFHQX1 \cpuregs_reg[10][27] (.CK (clk), .D (n_3833), .Q
       (\cpuregs[10] [27]));
  DFFHQX1 \cpuregs_reg[10][28] (.CK (clk), .D (n_3834), .Q
       (\cpuregs[10] [28]));
  DFFHQX1 \cpuregs_reg[10][29] (.CK (clk), .D (n_3832), .Q
       (\cpuregs[10] [29]));
  DFFHQX1 \cpuregs_reg[10][30] (.CK (clk), .D (n_3831), .Q
       (\cpuregs[10] [30]));
  DFFHQX1 \cpuregs_reg[10][31] (.CK (clk), .D (n_3830), .Q
       (\cpuregs[10] [31]));
  DFFHQX1 \cpuregs_reg[11][0] (.CK (clk), .D (n_3561), .Q
       (\cpuregs[11] [0]));
  DFFHQX1 \cpuregs_reg[11][1] (.CK (clk), .D (n_3829), .Q
       (\cpuregs[11] [1]));
  DFFHQX1 \cpuregs_reg[11][2] (.CK (clk), .D (n_3828), .Q
       (\cpuregs[11] [2]));
  DFFHQX1 \cpuregs_reg[11][3] (.CK (clk), .D (n_3827), .Q
       (\cpuregs[11] [3]));
  DFFHQX1 \cpuregs_reg[11][4] (.CK (clk), .D (n_3826), .Q
       (\cpuregs[11] [4]));
  DFFHQX1 \cpuregs_reg[11][5] (.CK (clk), .D (n_3825), .Q
       (\cpuregs[11] [5]));
  DFFHQX1 \cpuregs_reg[11][6] (.CK (clk), .D (n_3824), .Q
       (\cpuregs[11] [6]));
  DFFHQX1 \cpuregs_reg[11][7] (.CK (clk), .D (n_3823), .Q
       (\cpuregs[11] [7]));
  DFFHQX1 \cpuregs_reg[11][8] (.CK (clk), .D (n_4080), .Q
       (\cpuregs[11] [8]));
  DFFHQX1 \cpuregs_reg[11][9] (.CK (clk), .D (n_4082), .Q
       (\cpuregs[11] [9]));
  DFFHQX1 \cpuregs_reg[11][10] (.CK (clk), .D (n_4081), .Q
       (\cpuregs[11] [10]));
  DFFHQX1 \cpuregs_reg[11][11] (.CK (clk), .D (n_4079), .Q
       (\cpuregs[11] [11]));
  DFFHQX1 \cpuregs_reg[11][12] (.CK (clk), .D (n_4078), .Q
       (\cpuregs[11] [12]));
  DFFHQX1 \cpuregs_reg[11][13] (.CK (clk), .D (n_4077), .Q
       (\cpuregs[11] [13]));
  DFFHQX1 \cpuregs_reg[11][14] (.CK (clk), .D (n_4076), .Q
       (\cpuregs[11] [14]));
  DFFHQX1 \cpuregs_reg[11][15] (.CK (clk), .D (n_4075), .Q
       (\cpuregs[11] [15]));
  DFFHQX1 \cpuregs_reg[11][16] (.CK (clk), .D (n_4074), .Q
       (\cpuregs[11] [16]));
  DFFHQX1 \cpuregs_reg[11][17] (.CK (clk), .D (n_4073), .Q
       (\cpuregs[11] [17]));
  DFFHQX1 \cpuregs_reg[11][18] (.CK (clk), .D (n_4072), .Q
       (\cpuregs[11] [18]));
  DFFHQX1 \cpuregs_reg[11][19] (.CK (clk), .D (n_4071), .Q
       (\cpuregs[11] [19]));
  DFFHQX1 \cpuregs_reg[11][20] (.CK (clk), .D (n_4069), .Q
       (\cpuregs[11] [20]));
  DFFHQX1 \cpuregs_reg[11][21] (.CK (clk), .D (n_4068), .Q
       (\cpuregs[11] [21]));
  DFFHQX1 \cpuregs_reg[11][22] (.CK (clk), .D (n_4070), .Q
       (\cpuregs[11] [22]));
  DFFHQX1 \cpuregs_reg[11][23] (.CK (clk), .D (n_4067), .Q
       (\cpuregs[11] [23]));
  DFFHQX1 \cpuregs_reg[11][24] (.CK (clk), .D (n_4066), .Q
       (\cpuregs[11] [24]));
  DFFHQX1 \cpuregs_reg[11][25] (.CK (clk), .D (n_4065), .Q
       (\cpuregs[11] [25]));
  DFFHQX1 \cpuregs_reg[11][26] (.CK (clk), .D (n_4064), .Q
       (\cpuregs[11] [26]));
  DFFHQX1 \cpuregs_reg[11][27] (.CK (clk), .D (n_4063), .Q
       (\cpuregs[11] [27]));
  DFFHQX1 \cpuregs_reg[11][28] (.CK (clk), .D (n_4062), .Q
       (\cpuregs[11] [28]));
  DFFHQX1 \cpuregs_reg[11][29] (.CK (clk), .D (n_4061), .Q
       (\cpuregs[11] [29]));
  DFFHQX1 \cpuregs_reg[11][30] (.CK (clk), .D (n_4060), .Q
       (\cpuregs[11] [30]));
  DFFHQX1 \cpuregs_reg[11][31] (.CK (clk), .D (n_3997), .Q
       (\cpuregs[11] [31]));
  DFFHQX1 \cpuregs_reg[12][0] (.CK (clk), .D (n_3493), .Q
       (\cpuregs[12] [0]));
  DFFHQX1 \cpuregs_reg[12][1] (.CK (clk), .D (n_3698), .Q
       (\cpuregs[12] [1]));
  DFFHQX1 \cpuregs_reg[12][2] (.CK (clk), .D (n_3697), .Q
       (\cpuregs[12] [2]));
  DFFHQX1 \cpuregs_reg[12][3] (.CK (clk), .D (n_3696), .Q
       (\cpuregs[12] [3]));
  DFFHQX1 \cpuregs_reg[12][4] (.CK (clk), .D (n_3695), .Q
       (\cpuregs[12] [4]));
  DFFHQX1 \cpuregs_reg[12][5] (.CK (clk), .D (n_3694), .Q
       (\cpuregs[12] [5]));
  DFFHQX1 \cpuregs_reg[12][6] (.CK (clk), .D (n_3693), .Q
       (\cpuregs[12] [6]));
  DFFHQX1 \cpuregs_reg[12][7] (.CK (clk), .D (n_3690), .Q
       (\cpuregs[12] [7]));
  DFFHQX1 \cpuregs_reg[12][8] (.CK (clk), .D (n_3692), .Q
       (\cpuregs[12] [8]));
  DFFHQX1 \cpuregs_reg[12][9] (.CK (clk), .D (n_3691), .Q
       (\cpuregs[12] [9]));
  DFFHQX1 \cpuregs_reg[12][10] (.CK (clk), .D (n_3689), .Q
       (\cpuregs[12] [10]));
  DFFHQX1 \cpuregs_reg[12][11] (.CK (clk), .D (n_3688), .Q
       (\cpuregs[12] [11]));
  DFFHQX1 \cpuregs_reg[12][12] (.CK (clk), .D (n_3687), .Q
       (\cpuregs[12] [12]));
  DFFHQX1 \cpuregs_reg[12][13] (.CK (clk), .D (n_3686), .Q
       (\cpuregs[12] [13]));
  DFFHQX1 \cpuregs_reg[12][14] (.CK (clk), .D (n_3685), .Q
       (\cpuregs[12] [14]));
  DFFHQX1 \cpuregs_reg[12][15] (.CK (clk), .D (n_3684), .Q
       (\cpuregs[12] [15]));
  DFFHQX1 \cpuregs_reg[12][16] (.CK (clk), .D (n_3683), .Q
       (\cpuregs[12] [16]));
  DFFHQX1 \cpuregs_reg[12][17] (.CK (clk), .D (n_3682), .Q
       (\cpuregs[12] [17]));
  DFFHQX1 \cpuregs_reg[12][18] (.CK (clk), .D (n_3681), .Q
       (\cpuregs[12] [18]));
  DFFHQX1 \cpuregs_reg[12][19] (.CK (clk), .D (n_3680), .Q
       (\cpuregs[12] [19]));
  DFFHQX1 \cpuregs_reg[12][20] (.CK (clk), .D (n_3679), .Q
       (\cpuregs[12] [20]));
  DFFHQX1 \cpuregs_reg[12][21] (.CK (clk), .D (n_3678), .Q
       (\cpuregs[12] [21]));
  DFFHQX1 \cpuregs_reg[12][22] (.CK (clk), .D (n_3677), .Q
       (\cpuregs[12] [22]));
  DFFHQX1 \cpuregs_reg[12][23] (.CK (clk), .D (n_3676), .Q
       (\cpuregs[12] [23]));
  DFFHQX1 \cpuregs_reg[12][24] (.CK (clk), .D (n_3675), .Q
       (\cpuregs[12] [24]));
  DFFHQX1 \cpuregs_reg[12][25] (.CK (clk), .D (n_3674), .Q
       (\cpuregs[12] [25]));
  DFFHQX1 \cpuregs_reg[12][26] (.CK (clk), .D (n_3673), .Q
       (\cpuregs[12] [26]));
  DFFHQX1 \cpuregs_reg[12][27] (.CK (clk), .D (n_3672), .Q
       (\cpuregs[12] [27]));
  DFFHQX1 \cpuregs_reg[12][28] (.CK (clk), .D (n_3671), .Q
       (\cpuregs[12] [28]));
  DFFHQX1 \cpuregs_reg[12][29] (.CK (clk), .D (n_3670), .Q
       (\cpuregs[12] [29]));
  DFFHQX1 \cpuregs_reg[12][30] (.CK (clk), .D (n_3669), .Q
       (\cpuregs[12] [30]));
  DFFHQX1 \cpuregs_reg[12][31] (.CK (clk), .D (n_3668), .Q
       (\cpuregs[12] [31]));
  DFFHQX1 \cpuregs_reg[13][0] (.CK (clk), .D (n_3574), .Q
       (\cpuregs[13] [0]));
  DFFHQX1 \cpuregs_reg[13][1] (.CK (clk), .D (n_4059), .Q
       (\cpuregs[13] [1]));
  DFFHQX1 \cpuregs_reg[13][2] (.CK (clk), .D (n_4058), .Q
       (\cpuregs[13] [2]));
  DFFHQX1 \cpuregs_reg[13][3] (.CK (clk), .D (n_4057), .Q
       (\cpuregs[13] [3]));
  DFFHQX1 \cpuregs_reg[13][4] (.CK (clk), .D (n_4056), .Q
       (\cpuregs[13] [4]));
  DFFHQX1 \cpuregs_reg[13][5] (.CK (clk), .D (n_4055), .Q
       (\cpuregs[13] [5]));
  DFFHQX1 \cpuregs_reg[13][6] (.CK (clk), .D (n_4054), .Q
       (\cpuregs[13] [6]));
  DFFHQX1 \cpuregs_reg[13][7] (.CK (clk), .D (n_4053), .Q
       (\cpuregs[13] [7]));
  DFFHQX1 \cpuregs_reg[13][8] (.CK (clk), .D (n_4052), .Q
       (\cpuregs[13] [8]));
  DFFHQX1 \cpuregs_reg[13][9] (.CK (clk), .D (n_4051), .Q
       (\cpuregs[13] [9]));
  DFFHQX1 \cpuregs_reg[13][10] (.CK (clk), .D (n_4050), .Q
       (\cpuregs[13] [10]));
  DFFHQX1 \cpuregs_reg[13][11] (.CK (clk), .D (n_4049), .Q
       (\cpuregs[13] [11]));
  DFFHQX1 \cpuregs_reg[13][12] (.CK (clk), .D (n_4048), .Q
       (\cpuregs[13] [12]));
  DFFHQX1 \cpuregs_reg[13][13] (.CK (clk), .D (n_4047), .Q
       (\cpuregs[13] [13]));
  DFFHQX1 \cpuregs_reg[13][14] (.CK (clk), .D (n_4045), .Q
       (\cpuregs[13] [14]));
  DFFHQX1 \cpuregs_reg[13][15] (.CK (clk), .D (n_4046), .Q
       (\cpuregs[13] [15]));
  DFFHQX1 \cpuregs_reg[13][16] (.CK (clk), .D (n_4044), .Q
       (\cpuregs[13] [16]));
  DFFHQX1 \cpuregs_reg[13][17] (.CK (clk), .D (n_4043), .Q
       (\cpuregs[13] [17]));
  DFFHQX1 \cpuregs_reg[13][18] (.CK (clk), .D (n_4042), .Q
       (\cpuregs[13] [18]));
  DFFHQX1 \cpuregs_reg[13][19] (.CK (clk), .D (n_4041), .Q
       (\cpuregs[13] [19]));
  DFFHQX1 \cpuregs_reg[13][20] (.CK (clk), .D (n_4040), .Q
       (\cpuregs[13] [20]));
  DFFHQX1 \cpuregs_reg[13][21] (.CK (clk), .D (n_4039), .Q
       (\cpuregs[13] [21]));
  DFFHQX1 \cpuregs_reg[13][22] (.CK (clk), .D (n_4038), .Q
       (\cpuregs[13] [22]));
  DFFHQX1 \cpuregs_reg[13][23] (.CK (clk), .D (n_4037), .Q
       (\cpuregs[13] [23]));
  DFFHQX1 \cpuregs_reg[13][24] (.CK (clk), .D (n_4036), .Q
       (\cpuregs[13] [24]));
  DFFHQX1 \cpuregs_reg[13][25] (.CK (clk), .D (n_4282), .Q
       (\cpuregs[13] [25]));
  DFFHQX1 \cpuregs_reg[13][26] (.CK (clk), .D (n_4035), .Q
       (\cpuregs[13] [26]));
  DFFHQX1 \cpuregs_reg[13][27] (.CK (clk), .D (n_4034), .Q
       (\cpuregs[13] [27]));
  DFFHQX1 \cpuregs_reg[13][28] (.CK (clk), .D (n_4033), .Q
       (\cpuregs[13] [28]));
  DFFHQX1 \cpuregs_reg[13][29] (.CK (clk), .D (n_4032), .Q
       (\cpuregs[13] [29]));
  DFFHQX1 \cpuregs_reg[13][30] (.CK (clk), .D (n_4031), .Q
       (\cpuregs[13] [30]));
  DFFHQX1 \cpuregs_reg[13][31] (.CK (clk), .D (n_4030), .Q
       (\cpuregs[13] [31]));
  DFFHQX1 \cpuregs_reg[14][0] (.CK (clk), .D (n_3573), .Q
       (\cpuregs[14] [0]));
  DFFHQX1 \cpuregs_reg[14][1] (.CK (clk), .D (n_4029), .Q
       (\cpuregs[14] [1]));
  DFFHQX1 \cpuregs_reg[14][2] (.CK (clk), .D (n_4028), .Q
       (\cpuregs[14] [2]));
  DFFHQX1 \cpuregs_reg[14][3] (.CK (clk), .D (n_4027), .Q
       (\cpuregs[14] [3]));
  DFFHQX1 \cpuregs_reg[14][4] (.CK (clk), .D (n_4026), .Q
       (\cpuregs[14] [4]));
  DFFHQX1 \cpuregs_reg[14][5] (.CK (clk), .D (n_4025), .Q
       (\cpuregs[14] [5]));
  DFFHQX1 \cpuregs_reg[14][6] (.CK (clk), .D (n_4024), .Q
       (\cpuregs[14] [6]));
  DFFHQX1 \cpuregs_reg[14][7] (.CK (clk), .D (n_4023), .Q
       (\cpuregs[14] [7]));
  DFFHQX1 \cpuregs_reg[14][8] (.CK (clk), .D (n_4022), .Q
       (\cpuregs[14] [8]));
  DFFHQX1 \cpuregs_reg[14][9] (.CK (clk), .D (n_4021), .Q
       (\cpuregs[14] [9]));
  DFFHQX1 \cpuregs_reg[14][10] (.CK (clk), .D (n_4020), .Q
       (\cpuregs[14] [10]));
  DFFHQX1 \cpuregs_reg[14][11] (.CK (clk), .D (n_4019), .Q
       (\cpuregs[14] [11]));
  DFFHQX1 \cpuregs_reg[14][12] (.CK (clk), .D (n_4018), .Q
       (\cpuregs[14] [12]));
  DFFHQX1 \cpuregs_reg[14][13] (.CK (clk), .D (n_4017), .Q
       (\cpuregs[14] [13]));
  DFFHQX1 \cpuregs_reg[14][14] (.CK (clk), .D (n_4016), .Q
       (\cpuregs[14] [14]));
  DFFHQX1 \cpuregs_reg[14][15] (.CK (clk), .D (n_4015), .Q
       (\cpuregs[14] [15]));
  DFFHQX1 \cpuregs_reg[14][16] (.CK (clk), .D (n_4014), .Q
       (\cpuregs[14] [16]));
  DFFHQX1 \cpuregs_reg[14][17] (.CK (clk), .D (n_4013), .Q
       (\cpuregs[14] [17]));
  DFFHQX1 \cpuregs_reg[14][18] (.CK (clk), .D (n_4012), .Q
       (\cpuregs[14] [18]));
  DFFHQX1 \cpuregs_reg[14][19] (.CK (clk), .D (n_4011), .Q
       (\cpuregs[14] [19]));
  DFFHQX1 \cpuregs_reg[14][20] (.CK (clk), .D (n_4010), .Q
       (\cpuregs[14] [20]));
  DFFHQX1 \cpuregs_reg[14][21] (.CK (clk), .D (n_4009), .Q
       (\cpuregs[14] [21]));
  DFFHQX1 \cpuregs_reg[14][22] (.CK (clk), .D (n_4008), .Q
       (\cpuregs[14] [22]));
  DFFHQX1 \cpuregs_reg[14][23] (.CK (clk), .D (n_4007), .Q
       (\cpuregs[14] [23]));
  DFFHQX1 \cpuregs_reg[14][24] (.CK (clk), .D (n_4006), .Q
       (\cpuregs[14] [24]));
  DFFHQX1 \cpuregs_reg[14][25] (.CK (clk), .D (n_4005), .Q
       (\cpuregs[14] [25]));
  DFFHQX1 \cpuregs_reg[14][26] (.CK (clk), .D (n_4002), .Q
       (\cpuregs[14] [26]));
  DFFHQX1 \cpuregs_reg[14][27] (.CK (clk), .D (n_4004), .Q
       (\cpuregs[14] [27]));
  DFFHQX1 \cpuregs_reg[14][28] (.CK (clk), .D (n_4003), .Q
       (\cpuregs[14] [28]));
  DFFHQX1 \cpuregs_reg[14][29] (.CK (clk), .D (n_4001), .Q
       (\cpuregs[14] [29]));
  DFFHQX1 \cpuregs_reg[14][30] (.CK (clk), .D (n_4000), .Q
       (\cpuregs[14] [30]));
  DFFHQX1 \cpuregs_reg[14][31] (.CK (clk), .D (n_3999), .Q
       (\cpuregs[14] [31]));
  DFFHQX1 \cpuregs_reg[15][0] (.CK (clk), .D (n_3492), .Q
       (\cpuregs[15] [0]));
  DFFHQX1 \cpuregs_reg[15][1] (.CK (clk), .D (n_3666), .Q
       (\cpuregs[15] [1]));
  DFFHQX1 \cpuregs_reg[15][2] (.CK (clk), .D (n_3667), .Q
       (\cpuregs[15] [2]));
  DFFHQX1 \cpuregs_reg[15][3] (.CK (clk), .D (n_3665), .Q
       (\cpuregs[15] [3]));
  DFFHQX1 \cpuregs_reg[15][4] (.CK (clk), .D (n_3664), .Q
       (\cpuregs[15] [4]));
  DFFHQX1 \cpuregs_reg[15][5] (.CK (clk), .D (n_3663), .Q
       (\cpuregs[15] [5]));
  DFFHQX1 \cpuregs_reg[15][6] (.CK (clk), .D (n_3662), .Q
       (\cpuregs[15] [6]));
  DFFHQX1 \cpuregs_reg[15][7] (.CK (clk), .D (n_3661), .Q
       (\cpuregs[15] [7]));
  DFFHQX1 \cpuregs_reg[15][8] (.CK (clk), .D (n_3660), .Q
       (\cpuregs[15] [8]));
  DFFHQX1 \cpuregs_reg[15][9] (.CK (clk), .D (n_3659), .Q
       (\cpuregs[15] [9]));
  DFFHQX1 \cpuregs_reg[15][10] (.CK (clk), .D (n_3658), .Q
       (\cpuregs[15] [10]));
  DFFHQX1 \cpuregs_reg[15][11] (.CK (clk), .D (n_3657), .Q
       (\cpuregs[15] [11]));
  DFFHQX1 \cpuregs_reg[15][12] (.CK (clk), .D (n_3656), .Q
       (\cpuregs[15] [12]));
  DFFHQX1 \cpuregs_reg[15][13] (.CK (clk), .D (n_3655), .Q
       (\cpuregs[15] [13]));
  DFFHQX1 \cpuregs_reg[15][14] (.CK (clk), .D (n_3654), .Q
       (\cpuregs[15] [14]));
  DFFHQX1 \cpuregs_reg[15][15] (.CK (clk), .D (n_3653), .Q
       (\cpuregs[15] [15]));
  DFFHQX1 \cpuregs_reg[15][16] (.CK (clk), .D (n_3652), .Q
       (\cpuregs[15] [16]));
  DFFHQX1 \cpuregs_reg[15][17] (.CK (clk), .D (n_3651), .Q
       (\cpuregs[15] [17]));
  DFFHQX1 \cpuregs_reg[15][18] (.CK (clk), .D (n_3650), .Q
       (\cpuregs[15] [18]));
  DFFHQX1 \cpuregs_reg[15][19] (.CK (clk), .D (n_3649), .Q
       (\cpuregs[15] [19]));
  DFFHQX1 \cpuregs_reg[15][20] (.CK (clk), .D (n_3648), .Q
       (\cpuregs[15] [20]));
  DFFHQX1 \cpuregs_reg[15][21] (.CK (clk), .D (n_3647), .Q
       (\cpuregs[15] [21]));
  DFFHQX1 \cpuregs_reg[15][22] (.CK (clk), .D (n_3646), .Q
       (\cpuregs[15] [22]));
  DFFHQX1 \cpuregs_reg[15][23] (.CK (clk), .D (n_3645), .Q
       (\cpuregs[15] [23]));
  DFFHQX1 \cpuregs_reg[15][24] (.CK (clk), .D (n_3644), .Q
       (\cpuregs[15] [24]));
  DFFHQX1 \cpuregs_reg[15][25] (.CK (clk), .D (n_3643), .Q
       (\cpuregs[15] [25]));
  DFFHQX1 \cpuregs_reg[15][26] (.CK (clk), .D (n_3642), .Q
       (\cpuregs[15] [26]));
  DFFHQX1 \cpuregs_reg[15][27] (.CK (clk), .D (n_3641), .Q
       (\cpuregs[15] [27]));
  DFFHQX1 \cpuregs_reg[15][28] (.CK (clk), .D (n_3640), .Q
       (\cpuregs[15] [28]));
  DFFHQX1 \cpuregs_reg[15][29] (.CK (clk), .D (n_3639), .Q
       (\cpuregs[15] [29]));
  DFFHQX1 \cpuregs_reg[15][30] (.CK (clk), .D (n_3638), .Q
       (\cpuregs[15] [30]));
  DFFHQX1 \cpuregs_reg[15][31] (.CK (clk), .D (n_3637), .Q
       (\cpuregs[15] [31]));
  DFFHQX1 \cpuregs_reg[16][0] (.CK (clk), .D (n_3262), .Q
       (\cpuregs[16] [0]));
  DFFHQX1 \cpuregs_reg[16][1] (.CK (clk), .D (n_3326), .Q
       (\cpuregs[16] [1]));
  DFFHQX1 \cpuregs_reg[16][2] (.CK (clk), .D (n_3325), .Q
       (\cpuregs[16] [2]));
  DFFHQX1 \cpuregs_reg[16][3] (.CK (clk), .D (n_3324), .Q
       (\cpuregs[16] [3]));
  DFFHQX1 \cpuregs_reg[16][4] (.CK (clk), .D (n_3323), .Q
       (\cpuregs[16] [4]));
  DFFHQX1 \cpuregs_reg[16][5] (.CK (clk), .D (n_3322), .Q
       (\cpuregs[16] [5]));
  DFFHQX1 \cpuregs_reg[16][6] (.CK (clk), .D (n_3321), .Q
       (\cpuregs[16] [6]));
  DFFHQX1 \cpuregs_reg[16][7] (.CK (clk), .D (n_3320), .Q
       (\cpuregs[16] [7]));
  DFFHQX1 \cpuregs_reg[16][8] (.CK (clk), .D (n_3319), .Q
       (\cpuregs[16] [8]));
  DFFHQX1 \cpuregs_reg[16][9] (.CK (clk), .D (n_3318), .Q
       (\cpuregs[16] [9]));
  DFFHQX1 \cpuregs_reg[16][10] (.CK (clk), .D (n_3317), .Q
       (\cpuregs[16] [10]));
  DFFHQX1 \cpuregs_reg[16][11] (.CK (clk), .D (n_3316), .Q
       (\cpuregs[16] [11]));
  DFFHQX1 \cpuregs_reg[16][12] (.CK (clk), .D (n_3315), .Q
       (\cpuregs[16] [12]));
  DFFHQX1 \cpuregs_reg[16][13] (.CK (clk), .D (n_3314), .Q
       (\cpuregs[16] [13]));
  DFFHQX1 \cpuregs_reg[16][14] (.CK (clk), .D (n_3313), .Q
       (\cpuregs[16] [14]));
  DFFHQX1 \cpuregs_reg[16][15] (.CK (clk), .D (n_3312), .Q
       (\cpuregs[16] [15]));
  DFFHQX1 \cpuregs_reg[16][16] (.CK (clk), .D (n_3311), .Q
       (\cpuregs[16] [16]));
  DFFHQX1 \cpuregs_reg[16][17] (.CK (clk), .D (n_3310), .Q
       (\cpuregs[16] [17]));
  DFFHQX1 \cpuregs_reg[16][18] (.CK (clk), .D (n_3309), .Q
       (\cpuregs[16] [18]));
  DFFHQX1 \cpuregs_reg[16][19] (.CK (clk), .D (n_3307), .Q
       (\cpuregs[16] [19]));
  DFFHQX1 \cpuregs_reg[16][20] (.CK (clk), .D (n_3308), .Q
       (\cpuregs[16] [20]));
  DFFHQX1 \cpuregs_reg[16][21] (.CK (clk), .D (n_3306), .Q
       (\cpuregs[16] [21]));
  DFFHQX1 \cpuregs_reg[16][22] (.CK (clk), .D (n_3305), .Q
       (\cpuregs[16] [22]));
  DFFHQX1 \cpuregs_reg[16][23] (.CK (clk), .D (n_3304), .Q
       (\cpuregs[16] [23]));
  DFFHQX1 \cpuregs_reg[16][24] (.CK (clk), .D (n_3303), .Q
       (\cpuregs[16] [24]));
  DFFHQX1 \cpuregs_reg[16][25] (.CK (clk), .D (n_3300), .Q
       (\cpuregs[16] [25]));
  DFFHQX1 \cpuregs_reg[16][26] (.CK (clk), .D (n_3302), .Q
       (\cpuregs[16] [26]));
  DFFHQX1 \cpuregs_reg[16][27] (.CK (clk), .D (n_3301), .Q
       (\cpuregs[16] [27]));
  DFFHQX1 \cpuregs_reg[16][28] (.CK (clk), .D (n_3299), .Q
       (\cpuregs[16] [28]));
  DFFHQX1 \cpuregs_reg[16][29] (.CK (clk), .D (n_3298), .Q
       (\cpuregs[16] [29]));
  DFFHQX1 \cpuregs_reg[16][30] (.CK (clk), .D (n_3297), .Q
       (\cpuregs[16] [30]));
  DFFHQX1 \cpuregs_reg[16][31] (.CK (clk), .D (n_3296), .Q
       (\cpuregs[16] [31]));
  DFFHQX1 \cpuregs_reg[17][0] (.CK (clk), .D (n_3264), .Q
       (\cpuregs[17] [0]));
  DFFHQX1 \cpuregs_reg[17][1] (.CK (clk), .D (n_3390), .Q
       (\cpuregs[17] [1]));
  DFFHQX1 \cpuregs_reg[17][2] (.CK (clk), .D (n_3389), .Q
       (\cpuregs[17] [2]));
  DFFHQX1 \cpuregs_reg[17][3] (.CK (clk), .D (n_3388), .Q
       (\cpuregs[17] [3]));
  DFFHQX1 \cpuregs_reg[17][4] (.CK (clk), .D (n_3387), .Q
       (\cpuregs[17] [4]));
  DFFHQX1 \cpuregs_reg[17][5] (.CK (clk), .D (n_3386), .Q
       (\cpuregs[17] [5]));
  DFFHQX1 \cpuregs_reg[17][6] (.CK (clk), .D (n_3385), .Q
       (\cpuregs[17] [6]));
  DFFHQX1 \cpuregs_reg[17][7] (.CK (clk), .D (n_3384), .Q
       (\cpuregs[17] [7]));
  DFFHQX1 \cpuregs_reg[17][8] (.CK (clk), .D (n_3383), .Q
       (\cpuregs[17] [8]));
  DFFHQX1 \cpuregs_reg[17][9] (.CK (clk), .D (n_3382), .Q
       (\cpuregs[17] [9]));
  DFFHQX1 \cpuregs_reg[17][10] (.CK (clk), .D (n_3381), .Q
       (\cpuregs[17] [10]));
  DFFHQX1 \cpuregs_reg[17][11] (.CK (clk), .D (n_3380), .Q
       (\cpuregs[17] [11]));
  DFFHQX1 \cpuregs_reg[17][12] (.CK (clk), .D (n_3379), .Q
       (\cpuregs[17] [12]));
  DFFHQX1 \cpuregs_reg[17][13] (.CK (clk), .D (n_3378), .Q
       (\cpuregs[17] [13]));
  DFFHQX1 \cpuregs_reg[17][14] (.CK (clk), .D (n_3377), .Q
       (\cpuregs[17] [14]));
  DFFHQX1 \cpuregs_reg[17][15] (.CK (clk), .D (n_3376), .Q
       (\cpuregs[17] [15]));
  DFFHQX1 \cpuregs_reg[17][16] (.CK (clk), .D (n_3375), .Q
       (\cpuregs[17] [16]));
  DFFHQX1 \cpuregs_reg[17][17] (.CK (clk), .D (n_3374), .Q
       (\cpuregs[17] [17]));
  DFFHQX1 \cpuregs_reg[17][18] (.CK (clk), .D (n_3373), .Q
       (\cpuregs[17] [18]));
  DFFHQX1 \cpuregs_reg[17][19] (.CK (clk), .D (n_3371), .Q
       (\cpuregs[17] [19]));
  DFFHQX1 \cpuregs_reg[17][20] (.CK (clk), .D (n_3372), .Q
       (\cpuregs[17] [20]));
  DFFHQX1 \cpuregs_reg[17][21] (.CK (clk), .D (n_3370), .Q
       (\cpuregs[17] [21]));
  DFFHQX1 \cpuregs_reg[17][22] (.CK (clk), .D (n_3369), .Q
       (\cpuregs[17] [22]));
  DFFHQX1 \cpuregs_reg[17][23] (.CK (clk), .D (n_3367), .Q
       (\cpuregs[17] [23]));
  DFFHQX1 \cpuregs_reg[17][24] (.CK (clk), .D (n_3368), .Q
       (\cpuregs[17] [24]));
  DFFHQX1 \cpuregs_reg[17][25] (.CK (clk), .D (n_3366), .Q
       (\cpuregs[17] [25]));
  DFFHQX1 \cpuregs_reg[17][26] (.CK (clk), .D (n_3365), .Q
       (\cpuregs[17] [26]));
  DFFHQX1 \cpuregs_reg[17][27] (.CK (clk), .D (n_3364), .Q
       (\cpuregs[17] [27]));
  DFFHQX1 \cpuregs_reg[17][28] (.CK (clk), .D (n_3363), .Q
       (\cpuregs[17] [28]));
  DFFHQX1 \cpuregs_reg[17][29] (.CK (clk), .D (n_3362), .Q
       (\cpuregs[17] [29]));
  DFFHQX1 \cpuregs_reg[17][30] (.CK (clk), .D (n_3361), .Q
       (\cpuregs[17] [30]));
  DFFHQX1 \cpuregs_reg[17][31] (.CK (clk), .D (n_3360), .Q
       (\cpuregs[17] [31]));
  DFFHQX1 \cpuregs_reg[18][0] (.CK (clk), .D (n_3572), .Q
       (\cpuregs[18] [0]));
  DFFHQX1 \cpuregs_reg[18][1] (.CK (clk), .D (n_3996), .Q
       (\cpuregs[18] [1]));
  DFFHQX1 \cpuregs_reg[18][2] (.CK (clk), .D (n_3995), .Q
       (\cpuregs[18] [2]));
  DFFHQX1 \cpuregs_reg[18][3] (.CK (clk), .D (n_3994), .Q
       (\cpuregs[18] [3]));
  DFFHQX1 \cpuregs_reg[18][4] (.CK (clk), .D (n_3993), .Q
       (\cpuregs[18] [4]));
  DFFHQX1 \cpuregs_reg[18][5] (.CK (clk), .D (n_3992), .Q
       (\cpuregs[18] [5]));
  DFFHQX1 \cpuregs_reg[18][6] (.CK (clk), .D (n_3990), .Q
       (\cpuregs[18] [6]));
  DFFHQX1 \cpuregs_reg[18][7] (.CK (clk), .D (n_3989), .Q
       (\cpuregs[18] [7]));
  DFFHQX1 \cpuregs_reg[18][8] (.CK (clk), .D (n_3987), .Q
       (\cpuregs[18] [8]));
  DFFHQX1 \cpuregs_reg[18][9] (.CK (clk), .D (n_3986), .Q
       (\cpuregs[18] [9]));
  DFFHQX1 \cpuregs_reg[18][10] (.CK (clk), .D (n_3984), .Q
       (\cpuregs[18] [10]));
  DFFHQX1 \cpuregs_reg[18][11] (.CK (clk), .D (n_3983), .Q
       (\cpuregs[18] [11]));
  DFFHQX1 \cpuregs_reg[18][12] (.CK (clk), .D (n_3981), .Q
       (\cpuregs[18] [12]));
  DFFHQX1 \cpuregs_reg[18][13] (.CK (clk), .D (n_3979), .Q
       (\cpuregs[18] [13]));
  DFFHQX1 \cpuregs_reg[18][14] (.CK (clk), .D (n_3978), .Q
       (\cpuregs[18] [14]));
  DFFHQX1 \cpuregs_reg[18][15] (.CK (clk), .D (n_3976), .Q
       (\cpuregs[18] [15]));
  DFFHQX1 \cpuregs_reg[18][16] (.CK (clk), .D (n_3975), .Q
       (\cpuregs[18] [16]));
  DFFHQX1 \cpuregs_reg[18][17] (.CK (clk), .D (n_3973), .Q
       (\cpuregs[18] [17]));
  DFFHQX1 \cpuregs_reg[18][18] (.CK (clk), .D (n_3971), .Q
       (\cpuregs[18] [18]));
  DFFHQX1 \cpuregs_reg[18][19] (.CK (clk), .D (n_3970), .Q
       (\cpuregs[18] [19]));
  DFFHQX1 \cpuregs_reg[18][20] (.CK (clk), .D (n_3968), .Q
       (\cpuregs[18] [20]));
  DFFHQX1 \cpuregs_reg[18][21] (.CK (clk), .D (n_3967), .Q
       (\cpuregs[18] [21]));
  DFFHQX1 \cpuregs_reg[18][22] (.CK (clk), .D (n_3965), .Q
       (\cpuregs[18] [22]));
  DFFHQX1 \cpuregs_reg[18][23] (.CK (clk), .D (n_3964), .Q
       (\cpuregs[18] [23]));
  DFFHQX1 \cpuregs_reg[18][24] (.CK (clk), .D (n_4093), .Q
       (\cpuregs[18] [24]));
  DFFHQX1 \cpuregs_reg[18][25] (.CK (clk), .D (n_4094), .Q
       (\cpuregs[18] [25]));
  DFFHQX1 \cpuregs_reg[18][26] (.CK (clk), .D (n_4095), .Q
       (\cpuregs[18] [26]));
  DFFHQX1 \cpuregs_reg[18][27] (.CK (clk), .D (n_4098), .Q
       (\cpuregs[18] [27]));
  DFFHQX1 \cpuregs_reg[18][28] (.CK (clk), .D (n_4100), .Q
       (\cpuregs[18] [28]));
  DFFHQX1 \cpuregs_reg[18][29] (.CK (clk), .D (n_4101), .Q
       (\cpuregs[18] [29]));
  DFFHQX1 \cpuregs_reg[18][30] (.CK (clk), .D (n_4118), .Q
       (\cpuregs[18] [30]));
  DFFHQX1 \cpuregs_reg[18][31] (.CK (clk), .D (n_4119), .Q
       (\cpuregs[18] [31]));
  DFFHQX1 \cpuregs_reg[19][0] (.CK (clk), .D (n_3570), .Q
       (\cpuregs[19] [0]));
  DFFHQX1 \cpuregs_reg[19][1] (.CK (clk), .D (n_4121), .Q
       (\cpuregs[19] [1]));
  DFFHQX1 \cpuregs_reg[19][2] (.CK (clk), .D (n_4122), .Q
       (\cpuregs[19] [2]));
  DFFHQX1 \cpuregs_reg[19][3] (.CK (clk), .D (n_4123), .Q
       (\cpuregs[19] [3]));
  DFFHQX1 \cpuregs_reg[19][4] (.CK (clk), .D (n_4126), .Q
       (\cpuregs[19] [4]));
  DFFHQX1 \cpuregs_reg[19][5] (.CK (clk), .D (n_4127), .Q
       (\cpuregs[19] [5]));
  DFFHQX1 \cpuregs_reg[19][6] (.CK (clk), .D (n_4128), .Q
       (\cpuregs[19] [6]));
  DFFHQX1 \cpuregs_reg[19][7] (.CK (clk), .D (n_4129), .Q
       (\cpuregs[19] [7]));
  DFFHQX1 \cpuregs_reg[19][8] (.CK (clk), .D (n_4131), .Q
       (\cpuregs[19] [8]));
  DFFHQX1 \cpuregs_reg[19][9] (.CK (clk), .D (n_4133), .Q
       (\cpuregs[19] [9]));
  DFFHQX1 \cpuregs_reg[19][10] (.CK (clk), .D (n_4135), .Q
       (\cpuregs[19] [10]));
  DFFHQX1 \cpuregs_reg[19][11] (.CK (clk), .D (n_4136), .Q
       (\cpuregs[19] [11]));
  DFFHQX1 \cpuregs_reg[19][12] (.CK (clk), .D (n_4137), .Q
       (\cpuregs[19] [12]));
  DFFHQX1 \cpuregs_reg[19][13] (.CK (clk), .D (n_4138), .Q
       (\cpuregs[19] [13]));
  DFFHQX1 \cpuregs_reg[19][14] (.CK (clk), .D (n_4141), .Q
       (\cpuregs[19] [14]));
  DFFHQX1 \cpuregs_reg[19][15] (.CK (clk), .D (n_4143), .Q
       (\cpuregs[19] [15]));
  DFFHQX1 \cpuregs_reg[19][16] (.CK (clk), .D (n_4144), .Q
       (\cpuregs[19] [16]));
  DFFHQX1 \cpuregs_reg[19][17] (.CK (clk), .D (n_4145), .Q
       (\cpuregs[19] [17]));
  DFFHQX1 \cpuregs_reg[19][18] (.CK (clk), .D (n_4146), .Q
       (\cpuregs[19] [18]));
  DFFHQX1 \cpuregs_reg[19][19] (.CK (clk), .D (n_4148), .Q
       (\cpuregs[19] [19]));
  DFFHQX1 \cpuregs_reg[19][20] (.CK (clk), .D (n_4149), .Q
       (\cpuregs[19] [20]));
  DFFHQX1 \cpuregs_reg[19][21] (.CK (clk), .D (n_4150), .Q
       (\cpuregs[19] [21]));
  DFFHQX1 \cpuregs_reg[19][22] (.CK (clk), .D (n_4152), .Q
       (\cpuregs[19] [22]));
  DFFHQX1 \cpuregs_reg[19][23] (.CK (clk), .D (n_4154), .Q
       (\cpuregs[19] [23]));
  DFFHQX1 \cpuregs_reg[19][24] (.CK (clk), .D (n_4156), .Q
       (\cpuregs[19] [24]));
  DFFHQX1 \cpuregs_reg[19][25] (.CK (clk), .D (n_4158), .Q
       (\cpuregs[19] [25]));
  DFFHQX1 \cpuregs_reg[19][26] (.CK (clk), .D (n_4159), .Q
       (\cpuregs[19] [26]));
  DFFHQX1 \cpuregs_reg[19][27] (.CK (clk), .D (n_4160), .Q
       (\cpuregs[19] [27]));
  DFFHQX1 \cpuregs_reg[19][28] (.CK (clk), .D (n_4162), .Q
       (\cpuregs[19] [28]));
  DFFHQX1 \cpuregs_reg[19][29] (.CK (clk), .D (n_4163), .Q
       (\cpuregs[19] [29]));
  DFFHQX1 \cpuregs_reg[19][30] (.CK (clk), .D (n_4165), .Q
       (\cpuregs[19] [30]));
  DFFHQX1 \cpuregs_reg[19][31] (.CK (clk), .D (n_4167), .Q
       (\cpuregs[19] [31]));
  DFFHQX1 \cpuregs_reg[20][0] (.CK (clk), .D (n_3491), .Q
       (\cpuregs[20] [0]));
  DFFHQX1 \cpuregs_reg[20][1] (.CK (clk), .D (n_3636), .Q
       (\cpuregs[20] [1]));
  DFFHQX1 \cpuregs_reg[20][2] (.CK (clk), .D (n_3635), .Q
       (\cpuregs[20] [2]));
  DFFHQX1 \cpuregs_reg[20][3] (.CK (clk), .D (n_3634), .Q
       (\cpuregs[20] [3]));
  DFFHQX1 \cpuregs_reg[20][4] (.CK (clk), .D (n_3633), .Q
       (\cpuregs[20] [4]));
  DFFHQX1 \cpuregs_reg[20][5] (.CK (clk), .D (n_3632), .Q
       (\cpuregs[20] [5]));
  DFFHQX1 \cpuregs_reg[20][6] (.CK (clk), .D (n_3631), .Q
       (\cpuregs[20] [6]));
  DFFHQX1 \cpuregs_reg[20][7] (.CK (clk), .D (n_3630), .Q
       (\cpuregs[20] [7]));
  DFFHQX1 \cpuregs_reg[20][8] (.CK (clk), .D (n_3629), .Q
       (\cpuregs[20] [8]));
  DFFHQX1 \cpuregs_reg[20][9] (.CK (clk), .D (n_3628), .Q
       (\cpuregs[20] [9]));
  DFFHQX1 \cpuregs_reg[20][10] (.CK (clk), .D (n_3627), .Q
       (\cpuregs[20] [10]));
  DFFHQX1 \cpuregs_reg[20][11] (.CK (clk), .D (n_3626), .Q
       (\cpuregs[20] [11]));
  DFFHQX1 \cpuregs_reg[20][12] (.CK (clk), .D (n_3625), .Q
       (\cpuregs[20] [12]));
  DFFHQX1 \cpuregs_reg[20][13] (.CK (clk), .D (n_3624), .Q
       (\cpuregs[20] [13]));
  DFFHQX1 \cpuregs_reg[20][14] (.CK (clk), .D (n_3623), .Q
       (\cpuregs[20] [14]));
  DFFHQX1 \cpuregs_reg[20][15] (.CK (clk), .D (n_3622), .Q
       (\cpuregs[20] [15]));
  DFFHQX1 \cpuregs_reg[20][16] (.CK (clk), .D (n_3621), .Q
       (\cpuregs[20] [16]));
  DFFHQX1 \cpuregs_reg[20][17] (.CK (clk), .D (n_3620), .Q
       (\cpuregs[20] [17]));
  DFFHQX1 \cpuregs_reg[20][18] (.CK (clk), .D (n_3619), .Q
       (\cpuregs[20] [18]));
  DFFHQX1 \cpuregs_reg[20][19] (.CK (clk), .D (n_3618), .Q
       (\cpuregs[20] [19]));
  DFFHQX1 \cpuregs_reg[20][20] (.CK (clk), .D (n_3617), .Q
       (\cpuregs[20] [20]));
  DFFHQX1 \cpuregs_reg[20][21] (.CK (clk), .D (n_3616), .Q
       (\cpuregs[20] [21]));
  DFFHQX1 \cpuregs_reg[20][22] (.CK (clk), .D (n_3615), .Q
       (\cpuregs[20] [22]));
  DFFHQX1 \cpuregs_reg[20][23] (.CK (clk), .D (n_3614), .Q
       (\cpuregs[20] [23]));
  DFFHQX1 \cpuregs_reg[20][24] (.CK (clk), .D (n_3613), .Q
       (\cpuregs[20] [24]));
  DFFHQX1 \cpuregs_reg[20][25] (.CK (clk), .D (n_3612), .Q
       (\cpuregs[20] [25]));
  DFFHQX1 \cpuregs_reg[20][26] (.CK (clk), .D (n_3611), .Q
       (\cpuregs[20] [26]));
  DFFHQX1 \cpuregs_reg[20][27] (.CK (clk), .D (n_3610), .Q
       (\cpuregs[20] [27]));
  DFFHQX1 \cpuregs_reg[20][28] (.CK (clk), .D (n_3609), .Q
       (\cpuregs[20] [28]));
  DFFHQX1 \cpuregs_reg[20][29] (.CK (clk), .D (n_3608), .Q
       (\cpuregs[20] [29]));
  DFFHQX1 \cpuregs_reg[20][30] (.CK (clk), .D (n_3607), .Q
       (\cpuregs[20] [30]));
  DFFHQX1 \cpuregs_reg[20][31] (.CK (clk), .D (n_3606), .Q
       (\cpuregs[20] [31]));
  DFFHQX1 \cpuregs_reg[21][0] (.CK (clk), .D (n_3568), .Q
       (\cpuregs[21] [0]));
  DFFHQX1 \cpuregs_reg[21][1] (.CK (clk), .D (n_4185), .Q
       (\cpuregs[21] [1]));
  DFFHQX1 \cpuregs_reg[21][2] (.CK (clk), .D (n_4186), .Q
       (\cpuregs[21] [2]));
  DFFHQX1 \cpuregs_reg[21][3] (.CK (clk), .D (n_4187), .Q
       (\cpuregs[21] [3]));
  DFFHQX1 \cpuregs_reg[21][4] (.CK (clk), .D (n_4189), .Q
       (\cpuregs[21] [4]));
  DFFHQX1 \cpuregs_reg[21][5] (.CK (clk), .D (n_4190), .Q
       (\cpuregs[21] [5]));
  DFFHQX1 \cpuregs_reg[21][6] (.CK (clk), .D (n_4193), .Q
       (\cpuregs[21] [6]));
  DFFHQX1 \cpuregs_reg[21][7] (.CK (clk), .D (n_4195), .Q
       (\cpuregs[21] [7]));
  DFFHQX1 \cpuregs_reg[21][8] (.CK (clk), .D (n_4197), .Q
       (\cpuregs[21] [8]));
  DFFHQX1 \cpuregs_reg[21][9] (.CK (clk), .D (n_4198), .Q
       (\cpuregs[21] [9]));
  DFFHQX1 \cpuregs_reg[21][10] (.CK (clk), .D (n_4199), .Q
       (\cpuregs[21] [10]));
  DFFHQX1 \cpuregs_reg[21][11] (.CK (clk), .D (n_4201), .Q
       (\cpuregs[21] [11]));
  DFFHQX1 \cpuregs_reg[21][12] (.CK (clk), .D (n_4202), .Q
       (\cpuregs[21] [12]));
  DFFHQX1 \cpuregs_reg[21][13] (.CK (clk), .D (n_4204), .Q
       (\cpuregs[21] [13]));
  DFFHQX1 \cpuregs_reg[21][14] (.CK (clk), .D (n_4205), .Q
       (\cpuregs[21] [14]));
  DFFHQX1 \cpuregs_reg[21][15] (.CK (clk), .D (n_4207), .Q
       (\cpuregs[21] [15]));
  DFFHQX1 \cpuregs_reg[21][16] (.CK (clk), .D (n_4208), .Q
       (\cpuregs[21] [16]));
  DFFHQX1 \cpuregs_reg[21][17] (.CK (clk), .D (n_4210), .Q
       (\cpuregs[21] [17]));
  DFFHQX1 \cpuregs_reg[21][18] (.CK (clk), .D (n_4211), .Q
       (\cpuregs[21] [18]));
  DFFHQX1 \cpuregs_reg[21][19] (.CK (clk), .D (n_4212), .Q
       (\cpuregs[21] [19]));
  DFFHQX1 \cpuregs_reg[21][20] (.CK (clk), .D (n_4213), .Q
       (\cpuregs[21] [20]));
  DFFHQX1 \cpuregs_reg[21][21] (.CK (clk), .D (n_4215), .Q
       (\cpuregs[21] [21]));
  DFFHQX1 \cpuregs_reg[21][22] (.CK (clk), .D (n_4216), .Q
       (\cpuregs[21] [22]));
  DFFHQX1 \cpuregs_reg[21][23] (.CK (clk), .D (n_4219), .Q
       (\cpuregs[21] [23]));
  DFFHQX1 \cpuregs_reg[21][24] (.CK (clk), .D (n_4220), .Q
       (\cpuregs[21] [24]));
  DFFHQX1 \cpuregs_reg[21][25] (.CK (clk), .D (n_4221), .Q
       (\cpuregs[21] [25]));
  DFFHQX1 \cpuregs_reg[21][26] (.CK (clk), .D (n_4223), .Q
       (\cpuregs[21] [26]));
  DFFHQX1 \cpuregs_reg[21][27] (.CK (clk), .D (n_4224), .Q
       (\cpuregs[21] [27]));
  DFFHQX1 \cpuregs_reg[21][28] (.CK (clk), .D (n_4225), .Q
       (\cpuregs[21] [28]));
  DFFHQX1 \cpuregs_reg[21][29] (.CK (clk), .D (n_4228), .Q
       (\cpuregs[21] [29]));
  DFFHQX1 \cpuregs_reg[21][30] (.CK (clk), .D (n_4229), .Q
       (\cpuregs[21] [30]));
  DFFHQX1 \cpuregs_reg[21][31] (.CK (clk), .D (n_4231), .Q
       (\cpuregs[21] [31]));
  DFFHQX1 \cpuregs_reg[22][0] (.CK (clk), .D (n_3567), .Q
       (\cpuregs[22] [0]));
  DFFHQX1 \cpuregs_reg[22][1] (.CK (clk), .D (n_4233), .Q
       (\cpuregs[22] [1]));
  DFFHQX1 \cpuregs_reg[22][2] (.CK (clk), .D (n_4234), .Q
       (\cpuregs[22] [2]));
  DFFHQX1 \cpuregs_reg[22][3] (.CK (clk), .D (n_4235), .Q
       (\cpuregs[22] [3]));
  DFFHQX1 \cpuregs_reg[22][4] (.CK (clk), .D (n_4236), .Q
       (\cpuregs[22] [4]));
  DFFHQX1 \cpuregs_reg[22][5] (.CK (clk), .D (n_4237), .Q
       (\cpuregs[22] [5]));
  DFFHQX1 \cpuregs_reg[22][6] (.CK (clk), .D (n_4238), .Q
       (\cpuregs[22] [6]));
  DFFHQX1 \cpuregs_reg[22][7] (.CK (clk), .D (n_4239), .Q
       (\cpuregs[22] [7]));
  DFFHQX1 \cpuregs_reg[22][8] (.CK (clk), .D (n_4240), .Q
       (\cpuregs[22] [8]));
  DFFHQX1 \cpuregs_reg[22][9] (.CK (clk), .D (n_4241), .Q
       (\cpuregs[22] [9]));
  DFFHQX1 \cpuregs_reg[22][10] (.CK (clk), .D (n_4242), .Q
       (\cpuregs[22] [10]));
  DFFHQX1 \cpuregs_reg[22][11] (.CK (clk), .D (n_4243), .Q
       (\cpuregs[22] [11]));
  DFFHQX1 \cpuregs_reg[22][12] (.CK (clk), .D (n_4244), .Q
       (\cpuregs[22] [12]));
  DFFHQX1 \cpuregs_reg[22][13] (.CK (clk), .D (n_4245), .Q
       (\cpuregs[22] [13]));
  DFFHQX1 \cpuregs_reg[22][14] (.CK (clk), .D (n_4246), .Q
       (\cpuregs[22] [14]));
  DFFHQX1 \cpuregs_reg[22][15] (.CK (clk), .D (n_4247), .Q
       (\cpuregs[22] [15]));
  DFFHQX1 \cpuregs_reg[22][16] (.CK (clk), .D (n_4248), .Q
       (\cpuregs[22] [16]));
  DFFHQX1 \cpuregs_reg[22][17] (.CK (clk), .D (n_4249), .Q
       (\cpuregs[22] [17]));
  DFFHQX1 \cpuregs_reg[22][18] (.CK (clk), .D (n_4250), .Q
       (\cpuregs[22] [18]));
  DFFHQX1 \cpuregs_reg[22][19] (.CK (clk), .D (n_4251), .Q
       (\cpuregs[22] [19]));
  DFFHQX1 \cpuregs_reg[22][20] (.CK (clk), .D (n_4252), .Q
       (\cpuregs[22] [20]));
  DFFHQX1 \cpuregs_reg[22][21] (.CK (clk), .D (n_4253), .Q
       (\cpuregs[22] [21]));
  DFFHQX1 \cpuregs_reg[22][22] (.CK (clk), .D (n_4254), .Q
       (\cpuregs[22] [22]));
  DFFHQX1 \cpuregs_reg[22][23] (.CK (clk), .D (n_4255), .Q
       (\cpuregs[22] [23]));
  DFFHQX1 \cpuregs_reg[22][24] (.CK (clk), .D (n_4256), .Q
       (\cpuregs[22] [24]));
  DFFHQX1 \cpuregs_reg[22][25] (.CK (clk), .D (n_4257), .Q
       (\cpuregs[22] [25]));
  DFFHQX1 \cpuregs_reg[22][26] (.CK (clk), .D (n_4258), .Q
       (\cpuregs[22] [26]));
  DFFHQX1 \cpuregs_reg[22][27] (.CK (clk), .D (n_4259), .Q
       (\cpuregs[22] [27]));
  DFFHQX1 \cpuregs_reg[22][28] (.CK (clk), .D (n_4260), .Q
       (\cpuregs[22] [28]));
  DFFHQX1 \cpuregs_reg[22][29] (.CK (clk), .D (n_4261), .Q
       (\cpuregs[22] [29]));
  DFFHQX1 \cpuregs_reg[22][30] (.CK (clk), .D (n_4262), .Q
       (\cpuregs[22] [30]));
  DFFHQX1 \cpuregs_reg[22][31] (.CK (clk), .D (n_4263), .Q
       (\cpuregs[22] [31]));
  DFFHQX1 \cpuregs_reg[23][0] (.CK (clk), .D (n_3490), .Q
       (\cpuregs[23] [0]));
  DFFHQX1 \cpuregs_reg[23][1] (.CK (clk), .D (n_3605), .Q
       (\cpuregs[23] [1]));
  DFFHQX1 \cpuregs_reg[23][2] (.CK (clk), .D (n_3604), .Q
       (\cpuregs[23] [2]));
  DFFHQX1 \cpuregs_reg[23][3] (.CK (clk), .D (n_3603), .Q
       (\cpuregs[23] [3]));
  DFFHQX1 \cpuregs_reg[23][4] (.CK (clk), .D (n_3602), .Q
       (\cpuregs[23] [4]));
  DFFHQX1 \cpuregs_reg[23][5] (.CK (clk), .D (n_3601), .Q
       (\cpuregs[23] [5]));
  DFFHQX1 \cpuregs_reg[23][6] (.CK (clk), .D (n_3600), .Q
       (\cpuregs[23] [6]));
  DFFHQX1 \cpuregs_reg[23][7] (.CK (clk), .D (n_3599), .Q
       (\cpuregs[23] [7]));
  DFFHQX1 \cpuregs_reg[23][8] (.CK (clk), .D (n_3598), .Q
       (\cpuregs[23] [8]));
  DFFHQX1 \cpuregs_reg[23][9] (.CK (clk), .D (n_3597), .Q
       (\cpuregs[23] [9]));
  DFFHQX1 \cpuregs_reg[23][10] (.CK (clk), .D (n_3596), .Q
       (\cpuregs[23] [10]));
  DFFHQX1 \cpuregs_reg[23][11] (.CK (clk), .D (n_3595), .Q
       (\cpuregs[23] [11]));
  DFFHQX1 \cpuregs_reg[23][12] (.CK (clk), .D (n_3594), .Q
       (\cpuregs[23] [12]));
  DFFHQX1 \cpuregs_reg[23][13] (.CK (clk), .D (n_3593), .Q
       (\cpuregs[23] [13]));
  DFFHQX1 \cpuregs_reg[23][14] (.CK (clk), .D (n_3592), .Q
       (\cpuregs[23] [14]));
  DFFHQX1 \cpuregs_reg[23][15] (.CK (clk), .D (n_3591), .Q
       (\cpuregs[23] [15]));
  DFFHQX1 \cpuregs_reg[23][16] (.CK (clk), .D (n_3590), .Q
       (\cpuregs[23] [16]));
  DFFHQX1 \cpuregs_reg[23][17] (.CK (clk), .D (n_3589), .Q
       (\cpuregs[23] [17]));
  DFFHQX1 \cpuregs_reg[23][18] (.CK (clk), .D (n_3588), .Q
       (\cpuregs[23] [18]));
  DFFHQX1 \cpuregs_reg[23][19] (.CK (clk), .D (n_3587), .Q
       (\cpuregs[23] [19]));
  DFFHQX1 \cpuregs_reg[23][20] (.CK (clk), .D (n_3586), .Q
       (\cpuregs[23] [20]));
  DFFHQX1 \cpuregs_reg[23][21] (.CK (clk), .D (n_3585), .Q
       (\cpuregs[23] [21]));
  DFFHQX1 \cpuregs_reg[23][22] (.CK (clk), .D (n_3584), .Q
       (\cpuregs[23] [22]));
  DFFHQX1 \cpuregs_reg[23][23] (.CK (clk), .D (n_3583), .Q
       (\cpuregs[23] [23]));
  DFFHQX1 \cpuregs_reg[23][24] (.CK (clk), .D (n_3582), .Q
       (\cpuregs[23] [24]));
  DFFHQX1 \cpuregs_reg[23][25] (.CK (clk), .D (n_3581), .Q
       (\cpuregs[23] [25]));
  DFFHQX1 \cpuregs_reg[23][26] (.CK (clk), .D (n_3580), .Q
       (\cpuregs[23] [26]));
  DFFHQX1 \cpuregs_reg[23][27] (.CK (clk), .D (n_3579), .Q
       (\cpuregs[23] [27]));
  DFFHQX1 \cpuregs_reg[23][28] (.CK (clk), .D (n_3578), .Q
       (\cpuregs[23] [28]));
  DFFHQX1 \cpuregs_reg[23][29] (.CK (clk), .D (n_3577), .Q
       (\cpuregs[23] [29]));
  DFFHQX1 \cpuregs_reg[23][30] (.CK (clk), .D (n_3576), .Q
       (\cpuregs[23] [30]));
  DFFHQX1 \cpuregs_reg[23][31] (.CK (clk), .D (n_3575), .Q
       (\cpuregs[23] [31]));
  DFFHQX1 \cpuregs_reg[24][0] (.CK (clk), .D (n_3261), .Q
       (\cpuregs[24] [0]));
  DFFHQX1 \cpuregs_reg[24][1] (.CK (clk), .D (n_3295), .Q
       (\cpuregs[24] [1]));
  DFFHQX1 \cpuregs_reg[24][2] (.CK (clk), .D (n_3294), .Q
       (\cpuregs[24] [2]));
  DFFHQX1 \cpuregs_reg[24][3] (.CK (clk), .D (n_3293), .Q
       (\cpuregs[24] [3]));
  DFFHQX1 \cpuregs_reg[24][4] (.CK (clk), .D (n_3292), .Q
       (\cpuregs[24] [4]));
  DFFHQX1 \cpuregs_reg[24][5] (.CK (clk), .D (n_3291), .Q
       (\cpuregs[24] [5]));
  DFFHQX1 \cpuregs_reg[24][6] (.CK (clk), .D (n_3290), .Q
       (\cpuregs[24] [6]));
  DFFHQX1 \cpuregs_reg[24][7] (.CK (clk), .D (n_3289), .Q
       (\cpuregs[24] [7]));
  DFFHQX1 \cpuregs_reg[24][8] (.CK (clk), .D (n_3288), .Q
       (\cpuregs[24] [8]));
  DFFHQX1 \cpuregs_reg[24][9] (.CK (clk), .D (n_3287), .Q
       (\cpuregs[24] [9]));
  DFFHQX1 \cpuregs_reg[24][10] (.CK (clk), .D (n_3286), .Q
       (\cpuregs[24] [10]));
  DFFHQX1 \cpuregs_reg[24][11] (.CK (clk), .D (n_3285), .Q
       (\cpuregs[24] [11]));
  DFFHQX1 \cpuregs_reg[24][12] (.CK (clk), .D (n_3284), .Q
       (\cpuregs[24] [12]));
  DFFHQX1 \cpuregs_reg[24][13] (.CK (clk), .D (n_3283), .Q
       (\cpuregs[24] [13]));
  DFFHQX1 \cpuregs_reg[24][14] (.CK (clk), .D (n_3282), .Q
       (\cpuregs[24] [14]));
  DFFHQX1 \cpuregs_reg[24][15] (.CK (clk), .D (n_3281), .Q
       (\cpuregs[24] [15]));
  DFFHQX1 \cpuregs_reg[24][16] (.CK (clk), .D (n_3280), .Q
       (\cpuregs[24] [16]));
  DFFHQX1 \cpuregs_reg[24][17] (.CK (clk), .D (n_3279), .Q
       (\cpuregs[24] [17]));
  DFFHQX1 \cpuregs_reg[24][18] (.CK (clk), .D (n_3278), .Q
       (\cpuregs[24] [18]));
  DFFHQX1 \cpuregs_reg[24][19] (.CK (clk), .D (n_3277), .Q
       (\cpuregs[24] [19]));
  DFFHQX1 \cpuregs_reg[24][20] (.CK (clk), .D (n_3276), .Q
       (\cpuregs[24] [20]));
  DFFHQX1 \cpuregs_reg[24][21] (.CK (clk), .D (n_3265), .Q
       (\cpuregs[24] [21]));
  DFFHQX1 \cpuregs_reg[24][22] (.CK (clk), .D (n_3275), .Q
       (\cpuregs[24] [22]));
  DFFHQX1 \cpuregs_reg[24][23] (.CK (clk), .D (n_3274), .Q
       (\cpuregs[24] [23]));
  DFFHQX1 \cpuregs_reg[24][24] (.CK (clk), .D (n_3273), .Q
       (\cpuregs[24] [24]));
  DFFHQX1 \cpuregs_reg[24][25] (.CK (clk), .D (n_3272), .Q
       (\cpuregs[24] [25]));
  DFFHQX1 \cpuregs_reg[24][26] (.CK (clk), .D (n_3271), .Q
       (\cpuregs[24] [26]));
  DFFHQX1 \cpuregs_reg[24][27] (.CK (clk), .D (n_3270), .Q
       (\cpuregs[24] [27]));
  DFFHQX1 \cpuregs_reg[24][28] (.CK (clk), .D (n_3269), .Q
       (\cpuregs[24] [28]));
  DFFHQX1 \cpuregs_reg[24][29] (.CK (clk), .D (n_3268), .Q
       (\cpuregs[24] [29]));
  DFFHQX1 \cpuregs_reg[24][30] (.CK (clk), .D (n_3267), .Q
       (\cpuregs[24] [30]));
  DFFHQX1 \cpuregs_reg[24][31] (.CK (clk), .D (n_3266), .Q
       (\cpuregs[24] [31]));
  DFFHQX1 \cpuregs_reg[25][0] (.CK (clk), .D (n_3263), .Q
       (\cpuregs[25] [0]));
  DFFHQX1 \cpuregs_reg[25][1] (.CK (clk), .D (n_3355), .Q
       (\cpuregs[25] [1]));
  DFFHQX1 \cpuregs_reg[25][2] (.CK (clk), .D (n_3354), .Q
       (\cpuregs[25] [2]));
  DFFHQX1 \cpuregs_reg[25][3] (.CK (clk), .D (n_3353), .Q
       (\cpuregs[25] [3]));
  DFFHQX1 \cpuregs_reg[25][4] (.CK (clk), .D (n_3352), .Q
       (\cpuregs[25] [4]));
  DFFHQX1 \cpuregs_reg[25][5] (.CK (clk), .D (n_3351), .Q
       (\cpuregs[25] [5]));
  DFFHQX1 \cpuregs_reg[25][6] (.CK (clk), .D (n_3349), .Q
       (\cpuregs[25] [6]));
  DFFHQX1 \cpuregs_reg[25][7] (.CK (clk), .D (n_3348), .Q
       (\cpuregs[25] [7]));
  DFFHQX1 \cpuregs_reg[25][8] (.CK (clk), .D (n_3347), .Q
       (\cpuregs[25] [8]));
  DFFHQX1 \cpuregs_reg[25][9] (.CK (clk), .D (n_3346), .Q
       (\cpuregs[25] [9]));
  DFFHQX1 \cpuregs_reg[25][10] (.CK (clk), .D (n_3345), .Q
       (\cpuregs[25] [10]));
  DFFHQX1 \cpuregs_reg[25][11] (.CK (clk), .D (n_3344), .Q
       (\cpuregs[25] [11]));
  DFFHQX1 \cpuregs_reg[25][12] (.CK (clk), .D (n_3343), .Q
       (\cpuregs[25] [12]));
  DFFHQX1 \cpuregs_reg[25][13] (.CK (clk), .D (n_3350), .Q
       (\cpuregs[25] [13]));
  DFFHQX1 \cpuregs_reg[25][14] (.CK (clk), .D (n_3342), .Q
       (\cpuregs[25] [14]));
  DFFHQX1 \cpuregs_reg[25][15] (.CK (clk), .D (n_3341), .Q
       (\cpuregs[25] [15]));
  DFFHQX1 \cpuregs_reg[25][16] (.CK (clk), .D (n_3340), .Q
       (\cpuregs[25] [16]));
  DFFHQX1 \cpuregs_reg[25][17] (.CK (clk), .D (n_3339), .Q
       (\cpuregs[25] [17]));
  DFFHQX1 \cpuregs_reg[25][18] (.CK (clk), .D (n_3338), .Q
       (\cpuregs[25] [18]));
  DFFHQX1 \cpuregs_reg[25][19] (.CK (clk), .D (n_3337), .Q
       (\cpuregs[25] [19]));
  DFFHQX1 \cpuregs_reg[25][20] (.CK (clk), .D (n_3336), .Q
       (\cpuregs[25] [20]));
  DFFHQX1 \cpuregs_reg[25][21] (.CK (clk), .D (n_3356), .Q
       (\cpuregs[25] [21]));
  DFFHQX1 \cpuregs_reg[25][22] (.CK (clk), .D (n_3335), .Q
       (\cpuregs[25] [22]));
  DFFHQX1 \cpuregs_reg[25][23] (.CK (clk), .D (n_3334), .Q
       (\cpuregs[25] [23]));
  DFFHQX1 \cpuregs_reg[25][24] (.CK (clk), .D (n_3333), .Q
       (\cpuregs[25] [24]));
  DFFHQX1 \cpuregs_reg[25][25] (.CK (clk), .D (n_3357), .Q
       (\cpuregs[25] [25]));
  DFFHQX1 \cpuregs_reg[25][26] (.CK (clk), .D (n_3332), .Q
       (\cpuregs[25] [26]));
  DFFHQX1 \cpuregs_reg[25][27] (.CK (clk), .D (n_3331), .Q
       (\cpuregs[25] [27]));
  DFFHQX1 \cpuregs_reg[25][28] (.CK (clk), .D (n_3330), .Q
       (\cpuregs[25] [28]));
  DFFHQX1 \cpuregs_reg[25][29] (.CK (clk), .D (n_3358), .Q
       (\cpuregs[25] [29]));
  DFFHQX1 \cpuregs_reg[25][30] (.CK (clk), .D (n_3329), .Q
       (\cpuregs[25] [30]));
  DFFHQX1 \cpuregs_reg[25][31] (.CK (clk), .D (n_3328), .Q
       (\cpuregs[25] [31]));
  DFFHQX1 \cpuregs_reg[26][0] (.CK (clk), .D (n_3565), .Q
       (\cpuregs[26] [0]));
  DFFHQX1 \cpuregs_reg[26][1] (.CK (clk), .D (n_3947), .Q
       (\cpuregs[26] [1]));
  DFFHQX1 \cpuregs_reg[26][2] (.CK (clk), .D (n_3945), .Q
       (\cpuregs[26] [2]));
  DFFHQX1 \cpuregs_reg[26][3] (.CK (clk), .D (n_3944), .Q
       (\cpuregs[26] [3]));
  DFFHQX1 \cpuregs_reg[26][4] (.CK (clk), .D (n_3943), .Q
       (\cpuregs[26] [4]));
  DFFHQX1 \cpuregs_reg[26][5] (.CK (clk), .D (n_3942), .Q
       (\cpuregs[26] [5]));
  DFFHQX1 \cpuregs_reg[26][6] (.CK (clk), .D (n_3941), .Q
       (\cpuregs[26] [6]));
  DFFHQX1 \cpuregs_reg[26][7] (.CK (clk), .D (n_3940), .Q
       (\cpuregs[26] [7]));
  DFFHQX1 \cpuregs_reg[26][8] (.CK (clk), .D (n_3939), .Q
       (\cpuregs[26] [8]));
  DFFHQX1 \cpuregs_reg[26][9] (.CK (clk), .D (n_3938), .Q
       (\cpuregs[26] [9]));
  DFFHQX1 \cpuregs_reg[26][10] (.CK (clk), .D (n_3937), .Q
       (\cpuregs[26] [10]));
  DFFHQX1 \cpuregs_reg[26][11] (.CK (clk), .D (n_3935), .Q
       (\cpuregs[26] [11]));
  DFFHQX1 \cpuregs_reg[26][12] (.CK (clk), .D (n_3934), .Q
       (\cpuregs[26] [12]));
  DFFHQX1 \cpuregs_reg[26][13] (.CK (clk), .D (n_3933), .Q
       (\cpuregs[26] [13]));
  DFFHQX1 \cpuregs_reg[26][14] (.CK (clk), .D (n_3932), .Q
       (\cpuregs[26] [14]));
  DFFHQX1 \cpuregs_reg[26][15] (.CK (clk), .D (n_3929), .Q
       (\cpuregs[26] [15]));
  DFFHQX1 \cpuregs_reg[26][16] (.CK (clk), .D (n_3928), .Q
       (\cpuregs[26] [16]));
  DFFHQX1 \cpuregs_reg[26][17] (.CK (clk), .D (n_3927), .Q
       (\cpuregs[26] [17]));
  DFFHQX1 \cpuregs_reg[26][18] (.CK (clk), .D (n_3925), .Q
       (\cpuregs[26] [18]));
  DFFHQX1 \cpuregs_reg[26][19] (.CK (clk), .D (n_3923), .Q
       (\cpuregs[26] [19]));
  DFFHQX1 \cpuregs_reg[26][20] (.CK (clk), .D (n_3922), .Q
       (\cpuregs[26] [20]));
  DFFHQX1 \cpuregs_reg[26][21] (.CK (clk), .D (n_3921), .Q
       (\cpuregs[26] [21]));
  DFFHQX1 \cpuregs_reg[26][22] (.CK (clk), .D (n_3919), .Q
       (\cpuregs[26] [22]));
  DFFHQX1 \cpuregs_reg[26][23] (.CK (clk), .D (n_3918), .Q
       (\cpuregs[26] [23]));
  DFFHQX1 \cpuregs_reg[26][24] (.CK (clk), .D (n_3916), .Q
       (\cpuregs[26] [24]));
  DFFHQX1 \cpuregs_reg[26][25] (.CK (clk), .D (n_3914), .Q
       (\cpuregs[26] [25]));
  DFFHQX1 \cpuregs_reg[26][26] (.CK (clk), .D (n_3912), .Q
       (\cpuregs[26] [26]));
  DFFHQX1 \cpuregs_reg[26][27] (.CK (clk), .D (n_3911), .Q
       (\cpuregs[26] [27]));
  DFFHQX1 \cpuregs_reg[26][28] (.CK (clk), .D (n_3910), .Q
       (\cpuregs[26] [28]));
  DFFHQX1 \cpuregs_reg[26][29] (.CK (clk), .D (n_3908), .Q
       (\cpuregs[26] [29]));
  DFFHQX1 \cpuregs_reg[26][30] (.CK (clk), .D (n_3907), .Q
       (\cpuregs[26] [30]));
  DFFHQX1 \cpuregs_reg[26][31] (.CK (clk), .D (n_3905), .Q
       (\cpuregs[26] [31]));
  DFFHQX1 \cpuregs_reg[27][0] (.CK (clk), .D (n_3563), .Q
       (\cpuregs[27] [0]));
  DFFHQX1 \cpuregs_reg[27][1] (.CK (clk), .D (n_4191), .Q
       (\cpuregs[27] [1]));
  DFFHQX1 \cpuregs_reg[27][2] (.CK (clk), .D (n_3903), .Q
       (\cpuregs[27] [2]));
  DFFHQX1 \cpuregs_reg[27][3] (.CK (clk), .D (n_4182), .Q
       (\cpuregs[27] [3]));
  DFFHQX1 \cpuregs_reg[27][4] (.CK (clk), .D (n_3901), .Q
       (\cpuregs[27] [4]));
  DFFHQX1 \cpuregs_reg[27][5] (.CK (clk), .D (n_3900), .Q
       (\cpuregs[27] [5]));
  DFFHQX1 \cpuregs_reg[27][6] (.CK (clk), .D (n_3898), .Q
       (\cpuregs[27] [6]));
  DFFHQX1 \cpuregs_reg[27][7] (.CK (clk), .D (n_3897), .Q
       (\cpuregs[27] [7]));
  DFFHQX1 \cpuregs_reg[27][8] (.CK (clk), .D (n_3895), .Q
       (\cpuregs[27] [8]));
  DFFHQX1 \cpuregs_reg[27][9] (.CK (clk), .D (n_4173), .Q
       (\cpuregs[27] [9]));
  DFFHQX1 \cpuregs_reg[27][10] (.CK (clk), .D (n_3894), .Q
       (\cpuregs[27] [10]));
  DFFHQX1 \cpuregs_reg[27][11] (.CK (clk), .D (n_3892), .Q
       (\cpuregs[27] [11]));
  DFFHQX1 \cpuregs_reg[27][12] (.CK (clk), .D (n_3890), .Q
       (\cpuregs[27] [12]));
  DFFHQX1 \cpuregs_reg[27][13] (.CK (clk), .D (n_3889), .Q
       (\cpuregs[27] [13]));
  DFFHQX1 \cpuregs_reg[27][14] (.CK (clk), .D (n_3888), .Q
       (\cpuregs[27] [14]));
  DFFHQX1 \cpuregs_reg[27][15] (.CK (clk), .D (n_3861), .Q
       (\cpuregs[27] [15]));
  DFFHQX1 \cpuregs_reg[27][16] (.CK (clk), .D (n_3884), .Q
       (\cpuregs[27] [16]));
  DFFHQX1 \cpuregs_reg[27][17] (.CK (clk), .D (n_3955), .Q
       (\cpuregs[27] [17]));
  DFFHQX1 \cpuregs_reg[27][18] (.CK (clk), .D (n_3882), .Q
       (\cpuregs[27] [18]));
  DFFHQX1 \cpuregs_reg[27][19] (.CK (clk), .D (n_3881), .Q
       (\cpuregs[27] [19]));
  DFFHQX1 \cpuregs_reg[27][20] (.CK (clk), .D (n_3880), .Q
       (\cpuregs[27] [20]));
  DFFHQX1 \cpuregs_reg[27][21] (.CK (clk), .D (n_3878), .Q
       (\cpuregs[27] [21]));
  DFFHQX1 \cpuregs_reg[27][22] (.CK (clk), .D (n_3877), .Q
       (\cpuregs[27] [22]));
  DFFHQX1 \cpuregs_reg[27][23] (.CK (clk), .D (n_3876), .Q
       (\cpuregs[27] [23]));
  DFFHQX1 \cpuregs_reg[27][24] (.CK (clk), .D (n_3875), .Q
       (\cpuregs[27] [24]));
  DFFHQX1 \cpuregs_reg[27][25] (.CK (clk), .D (n_3873), .Q
       (\cpuregs[27] [25]));
  DFFHQX1 \cpuregs_reg[27][26] (.CK (clk), .D (n_3871), .Q
       (\cpuregs[27] [26]));
  DFFHQX1 \cpuregs_reg[27][27] (.CK (clk), .D (n_3870), .Q
       (\cpuregs[27] [27]));
  DFFHQX1 \cpuregs_reg[27][28] (.CK (clk), .D (n_3869), .Q
       (\cpuregs[27] [28]));
  DFFHQX1 \cpuregs_reg[27][29] (.CK (clk), .D (n_3868), .Q
       (\cpuregs[27] [29]));
  DFFHQX1 \cpuregs_reg[27][30] (.CK (clk), .D (n_3867), .Q
       (\cpuregs[27] [30]));
  DFFHQX1 \cpuregs_reg[27][31] (.CK (clk), .D (n_3866), .Q
       (\cpuregs[27] [31]));
  DFFHQX1 \cpuregs_reg[28][0] (.CK (clk), .D (n_3472), .Q
       (\cpuregs[28] [0]));
  DFFHQX1 \cpuregs_reg[28][1] (.CK (clk), .D (n_3560), .Q
       (\cpuregs[28] [1]));
  DFFHQX1 \cpuregs_reg[28][2] (.CK (clk), .D (n_3559), .Q
       (\cpuregs[28] [2]));
  DFFHQX1 \cpuregs_reg[28][3] (.CK (clk), .D (n_3558), .Q
       (\cpuregs[28] [3]));
  DFFHQX1 \cpuregs_reg[28][4] (.CK (clk), .D (n_3557), .Q
       (\cpuregs[28] [4]));
  DFFHQX1 \cpuregs_reg[28][5] (.CK (clk), .D (n_3556), .Q
       (\cpuregs[28] [5]));
  DFFHQX1 \cpuregs_reg[28][6] (.CK (clk), .D (n_3555), .Q
       (\cpuregs[28] [6]));
  DFFHQX1 \cpuregs_reg[28][7] (.CK (clk), .D (n_3554), .Q
       (\cpuregs[28] [7]));
  DFFHQX1 \cpuregs_reg[28][8] (.CK (clk), .D (n_3553), .Q
       (\cpuregs[28] [8]));
  DFFHQX1 \cpuregs_reg[28][9] (.CK (clk), .D (n_3552), .Q
       (\cpuregs[28] [9]));
  DFFHQX1 \cpuregs_reg[28][10] (.CK (clk), .D (n_3551), .Q
       (\cpuregs[28] [10]));
  DFFHQX1 \cpuregs_reg[28][11] (.CK (clk), .D (n_3550), .Q
       (\cpuregs[28] [11]));
  DFFHQX1 \cpuregs_reg[28][12] (.CK (clk), .D (n_3549), .Q
       (\cpuregs[28] [12]));
  DFFHQX1 \cpuregs_reg[28][13] (.CK (clk), .D (n_3548), .Q
       (\cpuregs[28] [13]));
  DFFHQX1 \cpuregs_reg[28][14] (.CK (clk), .D (n_3547), .Q
       (\cpuregs[28] [14]));
  DFFHQX1 \cpuregs_reg[28][15] (.CK (clk), .D (n_3546), .Q
       (\cpuregs[28] [15]));
  DFFHQX1 \cpuregs_reg[28][16] (.CK (clk), .D (n_3545), .Q
       (\cpuregs[28] [16]));
  DFFHQX1 \cpuregs_reg[28][17] (.CK (clk), .D (n_3544), .Q
       (\cpuregs[28] [17]));
  DFFHQX1 \cpuregs_reg[28][18] (.CK (clk), .D (n_3543), .Q
       (\cpuregs[28] [18]));
  DFFHQX1 \cpuregs_reg[28][19] (.CK (clk), .D (n_3542), .Q
       (\cpuregs[28] [19]));
  DFFHQX1 \cpuregs_reg[28][20] (.CK (clk), .D (n_3541), .Q
       (\cpuregs[28] [20]));
  DFFHQX1 \cpuregs_reg[28][21] (.CK (clk), .D (n_3540), .Q
       (\cpuregs[28] [21]));
  DFFHQX1 \cpuregs_reg[28][22] (.CK (clk), .D (n_3539), .Q
       (\cpuregs[28] [22]));
  DFFHQX1 \cpuregs_reg[28][23] (.CK (clk), .D (n_3538), .Q
       (\cpuregs[28] [23]));
  DFFHQX1 \cpuregs_reg[28][24] (.CK (clk), .D (n_3537), .Q
       (\cpuregs[28] [24]));
  DFFHQX1 \cpuregs_reg[28][25] (.CK (clk), .D (n_3536), .Q
       (\cpuregs[28] [25]));
  DFFHQX1 \cpuregs_reg[28][26] (.CK (clk), .D (n_3535), .Q
       (\cpuregs[28] [26]));
  DFFHQX1 \cpuregs_reg[28][27] (.CK (clk), .D (n_3534), .Q
       (\cpuregs[28] [27]));
  DFFHQX1 \cpuregs_reg[28][28] (.CK (clk), .D (n_3533), .Q
       (\cpuregs[28] [28]));
  DFFHQX1 \cpuregs_reg[28][29] (.CK (clk), .D (n_3532), .Q
       (\cpuregs[28] [29]));
  DFFHQX1 \cpuregs_reg[28][30] (.CK (clk), .D (n_3531), .Q
       (\cpuregs[28] [30]));
  DFFHQX1 \cpuregs_reg[28][31] (.CK (clk), .D (n_3530), .Q
       (\cpuregs[28] [31]));
  DFFHQX1 \cpuregs_reg[29][0] (.CK (clk), .D (n_3497), .Q
       (\cpuregs[29] [0]));
  DFFHQX1 \cpuregs_reg[29][1] (.CK (clk), .D (n_3791), .Q
       (\cpuregs[29] [1]));
  DFFHQX1 \cpuregs_reg[29][2] (.CK (clk), .D (n_3790), .Q
       (\cpuregs[29] [2]));
  DFFHQX1 \cpuregs_reg[29][3] (.CK (clk), .D (n_3789), .Q
       (\cpuregs[29] [3]));
  DFFHQX1 \cpuregs_reg[29][4] (.CK (clk), .D (n_3788), .Q
       (\cpuregs[29] [4]));
  DFFHQX1 \cpuregs_reg[29][5] (.CK (clk), .D (n_3787), .Q
       (\cpuregs[29] [5]));
  DFFHQX1 \cpuregs_reg[29][6] (.CK (clk), .D (n_3786), .Q
       (\cpuregs[29] [6]));
  DFFHQX1 \cpuregs_reg[29][7] (.CK (clk), .D (n_3785), .Q
       (\cpuregs[29] [7]));
  DFFHQX1 \cpuregs_reg[29][8] (.CK (clk), .D (n_3784), .Q
       (\cpuregs[29] [8]));
  DFFHQX1 \cpuregs_reg[29][9] (.CK (clk), .D (n_3783), .Q
       (\cpuregs[29] [9]));
  DFFHQX1 \cpuregs_reg[29][10] (.CK (clk), .D (n_3782), .Q
       (\cpuregs[29] [10]));
  DFFHQX1 \cpuregs_reg[29][11] (.CK (clk), .D (n_3781), .Q
       (\cpuregs[29] [11]));
  DFFHQX1 \cpuregs_reg[29][12] (.CK (clk), .D (n_3780), .Q
       (\cpuregs[29] [12]));
  DFFHQX1 \cpuregs_reg[29][13] (.CK (clk), .D (n_3779), .Q
       (\cpuregs[29] [13]));
  DFFHQX1 \cpuregs_reg[29][14] (.CK (clk), .D (n_3778), .Q
       (\cpuregs[29] [14]));
  DFFHQX1 \cpuregs_reg[29][15] (.CK (clk), .D (n_3777), .Q
       (\cpuregs[29] [15]));
  DFFHQX1 \cpuregs_reg[29][16] (.CK (clk), .D (n_3776), .Q
       (\cpuregs[29] [16]));
  DFFHQX1 \cpuregs_reg[29][17] (.CK (clk), .D (n_3775), .Q
       (\cpuregs[29] [17]));
  DFFHQX1 \cpuregs_reg[29][18] (.CK (clk), .D (n_3774), .Q
       (\cpuregs[29] [18]));
  DFFHQX1 \cpuregs_reg[29][19] (.CK (clk), .D (n_3773), .Q
       (\cpuregs[29] [19]));
  DFFHQX1 \cpuregs_reg[29][20] (.CK (clk), .D (n_3772), .Q
       (\cpuregs[29] [20]));
  DFFHQX1 \cpuregs_reg[29][21] (.CK (clk), .D (n_3771), .Q
       (\cpuregs[29] [21]));
  DFFHQX1 \cpuregs_reg[29][22] (.CK (clk), .D (n_3770), .Q
       (\cpuregs[29] [22]));
  DFFHQX1 \cpuregs_reg[29][23] (.CK (clk), .D (n_3769), .Q
       (\cpuregs[29] [23]));
  DFFHQX1 \cpuregs_reg[29][24] (.CK (clk), .D (n_3768), .Q
       (\cpuregs[29] [24]));
  DFFHQX1 \cpuregs_reg[29][25] (.CK (clk), .D (n_3767), .Q
       (\cpuregs[29] [25]));
  DFFHQX1 \cpuregs_reg[29][26] (.CK (clk), .D (n_3766), .Q
       (\cpuregs[29] [26]));
  DFFHQX1 \cpuregs_reg[29][27] (.CK (clk), .D (n_3765), .Q
       (\cpuregs[29] [27]));
  DFFHQX1 \cpuregs_reg[29][28] (.CK (clk), .D (n_3764), .Q
       (\cpuregs[29] [28]));
  DFFHQX1 \cpuregs_reg[29][29] (.CK (clk), .D (n_3763), .Q
       (\cpuregs[29] [29]));
  DFFHQX1 \cpuregs_reg[29][30] (.CK (clk), .D (n_3762), .Q
       (\cpuregs[29] [30]));
  DFFHQX1 \cpuregs_reg[29][31] (.CK (clk), .D (n_3761), .Q
       (\cpuregs[29] [31]));
  DFFHQX1 \cpuregs_reg[30][0] (.CK (clk), .D (n_3498), .Q
       (\cpuregs[30] [0]));
  DFFHQX1 \cpuregs_reg[30][1] (.CK (clk), .D (n_3822), .Q
       (\cpuregs[30] [1]));
  DFFHQX1 \cpuregs_reg[30][2] (.CK (clk), .D (n_3821), .Q
       (\cpuregs[30] [2]));
  DFFHQX1 \cpuregs_reg[30][3] (.CK (clk), .D (n_3820), .Q
       (\cpuregs[30] [3]));
  DFFHQX1 \cpuregs_reg[30][4] (.CK (clk), .D (n_3819), .Q
       (\cpuregs[30] [4]));
  DFFHQX1 \cpuregs_reg[30][5] (.CK (clk), .D (n_3818), .Q
       (\cpuregs[30] [5]));
  DFFHQX1 \cpuregs_reg[30][6] (.CK (clk), .D (n_3817), .Q
       (\cpuregs[30] [6]));
  DFFHQX1 \cpuregs_reg[30][7] (.CK (clk), .D (n_3816), .Q
       (\cpuregs[30] [7]));
  DFFHQX1 \cpuregs_reg[30][8] (.CK (clk), .D (n_3815), .Q
       (\cpuregs[30] [8]));
  DFFHQX1 \cpuregs_reg[30][9] (.CK (clk), .D (n_3809), .Q
       (\cpuregs[30] [9]));
  DFFHQX1 \cpuregs_reg[30][10] (.CK (clk), .D (n_3814), .Q
       (\cpuregs[30] [10]));
  DFFHQX1 \cpuregs_reg[30][11] (.CK (clk), .D (n_3813), .Q
       (\cpuregs[30] [11]));
  DFFHQX1 \cpuregs_reg[30][12] (.CK (clk), .D (n_3812), .Q
       (\cpuregs[30] [12]));
  DFFHQX1 \cpuregs_reg[30][13] (.CK (clk), .D (n_3811), .Q
       (\cpuregs[30] [13]));
  DFFHQX1 \cpuregs_reg[30][14] (.CK (clk), .D (n_3810), .Q
       (\cpuregs[30] [14]));
  DFFHQX1 \cpuregs_reg[30][15] (.CK (clk), .D (n_3808), .Q
       (\cpuregs[30] [15]));
  DFFHQX1 \cpuregs_reg[30][16] (.CK (clk), .D (n_3807), .Q
       (\cpuregs[30] [16]));
  DFFHQX1 \cpuregs_reg[30][17] (.CK (clk), .D (n_3806), .Q
       (\cpuregs[30] [17]));
  DFFHQX1 \cpuregs_reg[30][18] (.CK (clk), .D (n_3805), .Q
       (\cpuregs[30] [18]));
  DFFHQX1 \cpuregs_reg[30][19] (.CK (clk), .D (n_3804), .Q
       (\cpuregs[30] [19]));
  DFFHQX1 \cpuregs_reg[30][20] (.CK (clk), .D (n_3803), .Q
       (\cpuregs[30] [20]));
  DFFHQX1 \cpuregs_reg[30][21] (.CK (clk), .D (n_3802), .Q
       (\cpuregs[30] [21]));
  DFFHQX1 \cpuregs_reg[30][22] (.CK (clk), .D (n_3799), .Q
       (\cpuregs[30] [22]));
  DFFHQX1 \cpuregs_reg[30][23] (.CK (clk), .D (n_3801), .Q
       (\cpuregs[30] [23]));
  DFFHQX1 \cpuregs_reg[30][24] (.CK (clk), .D (n_3800), .Q
       (\cpuregs[30] [24]));
  DFFHQX1 \cpuregs_reg[30][25] (.CK (clk), .D (n_3797), .Q
       (\cpuregs[30] [25]));
  DFFHQX1 \cpuregs_reg[30][26] (.CK (clk), .D (n_3798), .Q
       (\cpuregs[30] [26]));
  DFFHQX1 \cpuregs_reg[30][27] (.CK (clk), .D (n_3796), .Q
       (\cpuregs[30] [27]));
  DFFHQX1 \cpuregs_reg[30][28] (.CK (clk), .D (n_3795), .Q
       (\cpuregs[30] [28]));
  DFFHQX1 \cpuregs_reg[30][29] (.CK (clk), .D (n_3793), .Q
       (\cpuregs[30] [29]));
  DFFHQX1 \cpuregs_reg[30][30] (.CK (clk), .D (n_3794), .Q
       (\cpuregs[30] [30]));
  DFFHQX1 \cpuregs_reg[30][31] (.CK (clk), .D (n_3792), .Q
       (\cpuregs[30] [31]));
  DFFHQX1 \cpuregs_reg[31][0] (.CK (clk), .D (n_3471), .Q
       (\cpuregs[31] [0]));
  DFFHQX1 \cpuregs_reg[31][1] (.CK (clk), .D (n_3529), .Q
       (\cpuregs[31] [1]));
  DFFHQX1 \cpuregs_reg[31][2] (.CK (clk), .D (n_3528), .Q
       (\cpuregs[31] [2]));
  DFFHQX1 \cpuregs_reg[31][3] (.CK (clk), .D (n_3527), .Q
       (\cpuregs[31] [3]));
  DFFHQX1 \cpuregs_reg[31][4] (.CK (clk), .D (n_3526), .Q
       (\cpuregs[31] [4]));
  DFFHQX1 \cpuregs_reg[31][5] (.CK (clk), .D (n_3525), .Q
       (\cpuregs[31] [5]));
  DFFHQX1 \cpuregs_reg[31][6] (.CK (clk), .D (n_3524), .Q
       (\cpuregs[31] [6]));
  DFFHQX1 \cpuregs_reg[31][7] (.CK (clk), .D (n_3523), .Q
       (\cpuregs[31] [7]));
  DFFHQX1 \cpuregs_reg[31][8] (.CK (clk), .D (n_3522), .Q
       (\cpuregs[31] [8]));
  DFFHQX1 \cpuregs_reg[31][9] (.CK (clk), .D (n_3521), .Q
       (\cpuregs[31] [9]));
  DFFHQX1 \cpuregs_reg[31][10] (.CK (clk), .D (n_3520), .Q
       (\cpuregs[31] [10]));
  DFFHQX1 \cpuregs_reg[31][11] (.CK (clk), .D (n_3519), .Q
       (\cpuregs[31] [11]));
  DFFHQX1 \cpuregs_reg[31][12] (.CK (clk), .D (n_3518), .Q
       (\cpuregs[31] [12]));
  DFFHQX1 \cpuregs_reg[31][13] (.CK (clk), .D (n_3517), .Q
       (\cpuregs[31] [13]));
  DFFHQX1 \cpuregs_reg[31][14] (.CK (clk), .D (n_3516), .Q
       (\cpuregs[31] [14]));
  DFFHQX1 \cpuregs_reg[31][15] (.CK (clk), .D (n_3515), .Q
       (\cpuregs[31] [15]));
  DFFHQX1 \cpuregs_reg[31][16] (.CK (clk), .D (n_3514), .Q
       (\cpuregs[31] [16]));
  DFFHQX1 \cpuregs_reg[31][17] (.CK (clk), .D (n_3513), .Q
       (\cpuregs[31] [17]));
  DFFHQX1 \cpuregs_reg[31][18] (.CK (clk), .D (n_3512), .Q
       (\cpuregs[31] [18]));
  DFFHQX1 \cpuregs_reg[31][19] (.CK (clk), .D (n_3511), .Q
       (\cpuregs[31] [19]));
  DFFHQX1 \cpuregs_reg[31][20] (.CK (clk), .D (n_3509), .Q
       (\cpuregs[31] [20]));
  DFFHQX1 \cpuregs_reg[31][21] (.CK (clk), .D (n_3510), .Q
       (\cpuregs[31] [21]));
  DFFHQX1 \cpuregs_reg[31][22] (.CK (clk), .D (n_3508), .Q
       (\cpuregs[31] [22]));
  DFFHQX1 \cpuregs_reg[31][23] (.CK (clk), .D (n_3507), .Q
       (\cpuregs[31] [23]));
  DFFHQX1 \cpuregs_reg[31][24] (.CK (clk), .D (n_3506), .Q
       (\cpuregs[31] [24]));
  DFFHQX1 \cpuregs_reg[31][25] (.CK (clk), .D (n_3505), .Q
       (\cpuregs[31] [25]));
  DFFHQX1 \cpuregs_reg[31][26] (.CK (clk), .D (n_3504), .Q
       (\cpuregs[31] [26]));
  DFFHQX1 \cpuregs_reg[31][27] (.CK (clk), .D (n_3503), .Q
       (\cpuregs[31] [27]));
  DFFHQX1 \cpuregs_reg[31][28] (.CK (clk), .D (n_3502), .Q
       (\cpuregs[31] [28]));
  DFFHQX1 \cpuregs_reg[31][29] (.CK (clk), .D (n_3500), .Q
       (\cpuregs[31] [29]));
  DFFHQX1 \cpuregs_reg[31][30] (.CK (clk), .D (n_3501), .Q
       (\cpuregs[31] [30]));
  DFFHQX1 \cpuregs_reg[31][31] (.CK (clk), .D (n_3499), .Q
       (\cpuregs[31] [31]));
  DFFHQX1 \decoded_imm_j_reg[1] (.CK (clk), .D (n_2339), .Q
       (decoded_imm_j[1]));
  DFFHQX1 \decoded_imm_j_reg[2] (.CK (clk), .D (n_2395), .Q
       (decoded_imm_j[2]));
  DFFHQX1 \decoded_imm_j_reg[3] (.CK (clk), .D (n_2476), .Q
       (decoded_imm_j[3]));
  DFFHQX1 \decoded_imm_j_reg[4] (.CK (clk), .D (n_2372), .Q
       (decoded_imm_j[4]));
  DFFHQX1 \decoded_imm_j_reg[5] (.CK (clk), .D (n_2417), .Q
       (decoded_imm_j[5]));
  DFFHQX1 \decoded_imm_j_reg[6] (.CK (clk), .D (n_2397), .Q
       (decoded_imm_j[6]));
  DFFHQX1 \decoded_imm_j_reg[7] (.CK (clk), .D (n_2416), .Q
       (decoded_imm_j[7]));
  DFFHQX1 \decoded_imm_j_reg[8] (.CK (clk), .D (n_2354), .Q
       (decoded_imm_j[8]));
  DFFHQX1 \decoded_imm_j_reg[9] (.CK (clk), .D (n_2366), .Q
       (decoded_imm_j[9]));
  DFFHQX1 \decoded_imm_j_reg[10] (.CK (clk), .D (n_2383), .Q
       (decoded_imm_j[10]));
  DFFHQX1 \decoded_imm_j_reg[11] (.CK (clk), .D (n_2398), .Q
       (decoded_imm_j[11]));
  DFFHQX1 \decoded_imm_j_reg[12] (.CK (clk), .D (n_2345), .Q
       (decoded_imm_j[12]));
  DFFHQX1 \decoded_imm_j_reg[13] (.CK (clk), .D (n_2475), .Q
       (decoded_imm_j[13]));
  DFFHQX1 \decoded_imm_j_reg[14] (.CK (clk), .D (n_2477), .Q
       (decoded_imm_j[14]));
  DFFHQX1 \decoded_imm_j_reg[15] (.CK (clk), .D (n_2478), .Q
       (decoded_imm_j[15]));
  DFFHQX1 \decoded_imm_j_reg[16] (.CK (clk), .D (n_2411), .Q
       (decoded_imm_j[16]));
  DFFHQX1 \decoded_imm_j_reg[17] (.CK (clk), .D (n_2412), .Q
       (decoded_imm_j[17]));
  DFFHQX1 \decoded_imm_j_reg[18] (.CK (clk), .D (n_2404), .Q
       (decoded_imm_j[18]));
  DFFHQX1 \decoded_imm_j_reg[19] (.CK (clk), .D (n_2387), .Q
       (decoded_imm_j[19]));
  DFFHQX1 \decoded_imm_j_reg[20] (.CK (clk), .D (n_2394), .Q
       (decoded_imm_j[20]));
  DFFHQX1 \decoded_imm_reg[1] (.CK (clk), .D (n_2276), .Q
       (decoded_imm[1]));
  DFFHQX1 \decoded_imm_reg[2] (.CK (clk), .D (n_2275), .Q
       (decoded_imm[2]));
  DFFHQX1 \decoded_imm_reg[3] (.CK (clk), .D (n_2274), .Q
       (decoded_imm[3]));
  DFFHQX1 \decoded_imm_reg[4] (.CK (clk), .D (n_2277), .Q
       (decoded_imm[4]));
  DFFHQX1 \decoded_imm_reg[5] (.CK (clk), .D (n_2228), .Q
       (decoded_imm[5]));
  DFFHQX1 \decoded_imm_reg[6] (.CK (clk), .D (n_2224), .Q
       (decoded_imm[6]));
  DFFHQX1 \decoded_imm_reg[7] (.CK (clk), .D (n_2223), .Q
       (decoded_imm[7]));
  DFFHQX1 \decoded_imm_reg[8] (.CK (clk), .D (n_2229), .Q
       (decoded_imm[8]));
  DFFHQX1 \decoded_imm_reg[9] (.CK (clk), .D (n_2258), .Q
       (decoded_imm[9]));
  DFFHQX1 \decoded_imm_reg[10] (.CK (clk), .D (n_2259), .Q
       (decoded_imm[10]));
  DFFHQX1 \decoded_imm_reg[11] (.CK (clk), .D (n_2384), .Q
       (decoded_imm[11]));
  DFFHQX1 \decoded_imm_reg[12] (.CK (clk), .D (n_2296), .Q
       (decoded_imm[12]));
  DFFHQX1 \decoded_imm_reg[13] (.CK (clk), .D (n_2298), .Q
       (decoded_imm[13]));
  DFFHQX1 \decoded_imm_reg[14] (.CK (clk), .D (n_2299), .Q
       (decoded_imm[14]));
  DFFHQX1 \decoded_imm_reg[15] (.CK (clk), .D (n_2300), .Q
       (decoded_imm[15]));
  DFFHQX1 \decoded_imm_reg[16] (.CK (clk), .D (n_2301), .Q
       (decoded_imm[16]));
  DFFHQX1 \decoded_imm_reg[17] (.CK (clk), .D (n_2302), .Q
       (decoded_imm[17]));
  DFFHQX1 \decoded_imm_reg[18] (.CK (clk), .D (n_2303), .Q
       (decoded_imm[18]));
  DFFHQX1 \decoded_imm_reg[19] (.CK (clk), .D (n_2304), .Q
       (decoded_imm[19]));
  DFFHQX1 \decoded_imm_reg[20] (.CK (clk), .D (n_2410), .Q
       (decoded_imm[20]));
  DFFHQX1 \decoded_imm_reg[21] (.CK (clk), .D (n_2403), .Q
       (decoded_imm[21]));
  DFFHQX1 \decoded_imm_reg[22] (.CK (clk), .D (n_2402), .Q
       (decoded_imm[22]));
  DFFHQX1 \decoded_imm_reg[23] (.CK (clk), .D (n_2400), .Q
       (decoded_imm[23]));
  DFFHQX1 \decoded_imm_reg[24] (.CK (clk), .D (n_2409), .Q
       (decoded_imm[24]));
  DFFHQX1 \decoded_imm_reg[25] (.CK (clk), .D (n_2408), .Q
       (decoded_imm[25]));
  DFFHQX1 \decoded_imm_reg[26] (.CK (clk), .D (n_2407), .Q
       (decoded_imm[26]));
  DFFHQX1 \decoded_imm_reg[27] (.CK (clk), .D (n_2399), .Q
       (decoded_imm[27]));
  DFFHQX1 \decoded_imm_reg[28] (.CK (clk), .D (n_2406), .Q
       (decoded_imm[28]));
  DFFHQX1 \decoded_imm_reg[29] (.CK (clk), .D (n_2405), .Q
       (decoded_imm[29]));
  DFFHQX1 \decoded_imm_reg[30] (.CK (clk), .D (n_2401), .Q
       (decoded_imm[30]));
  DFFHQX1 \decoded_imm_reg[31] (.CK (clk), .D (n_2396), .Q
       (decoded_imm[31]));
  DFFHQX1 \decoded_rd_reg[0] (.CK (clk), .D (n_5091), .Q
       (decoded_rd[0]));
  DFFHQX1 \decoded_rd_reg[1] (.CK (clk), .D (n_5046), .Q
       (decoded_rd[1]));
  DFFHQX1 \decoded_rd_reg[2] (.CK (clk), .D (n_5032), .Q
       (decoded_rd[2]));
  DFFHQX1 \decoded_rd_reg[3] (.CK (clk), .D (n_5054), .Q
       (decoded_rd[3]));
  DFFHQX1 \decoded_rd_reg[4] (.CK (clk), .D (n_4976), .Q
       (decoded_rd[4]));
  DFFHQX1 \decoded_rs1_reg[0] (.CK (clk), .D (n_4899), .Q
       (decoded_rs1[0]));
  DFFHQX1 \decoded_rs1_reg[1] (.CK (clk), .D (n_4974), .Q
       (decoded_rs1[1]));
  DFFHQX1 \decoded_rs1_reg[2] (.CK (clk), .D (n_4907), .Q
       (decoded_rs1[2]));
  DFFHQX1 \decoded_rs1_reg[3] (.CK (clk), .D (n_4910), .Q
       (decoded_rs1[3]));
  DFFHQX1 \decoded_rs2_reg[1] (.CK (clk), .D (n_4849), .Q
       (decoded_rs2[1]));
  DFFHQX1 decoder_trigger_reg(.CK (clk), .D (n_5528), .Q
       (decoder_trigger));
  DFFHQX1 \genblk1.pcpi_mul_active_reg[0] (.CK (clk), .D (n_1310), .Q
       (\genblk1.pcpi_mul_active [0]));
  DFFHQX1 \genblk1.pcpi_mul_active_reg[1] (.CK (clk), .D (n_807), .Q
       (pcpi_mul_wr));
  MDFFHQX4 \genblk1.pcpi_mul_rs1_reg[0] (.CK (clk), .D0 (reg_op1[0]),
       .D1 (\genblk1.pcpi_mul_rs1 [0]), .S0 (n_672), .Q
       (\genblk1.pcpi_mul_rs1 [0]));
  MDFFHQX4 \genblk1.pcpi_mul_rs2_reg[1] (.CK (clk), .D0
       (\reg_op2[1]_9670 ), .D1 (\genblk1.pcpi_mul_rs2 [1]), .S0
       (n_672), .Q (\genblk1.pcpi_mul_rs2 [1]));
  DFFHQX1 \genblk1.pcpi_mul_rs2_reg[2] (.CK (clk), .D (n_1664), .Q
       (\genblk1.pcpi_mul_rs2 [2]));
  MDFFHQX4 \genblk1.pcpi_mul_rs2_reg[3] (.CK (clk), .D0
       (\reg_op2[3]_9672 ), .D1 (\genblk1.pcpi_mul_rs2 [3]), .S0
       (n_672), .Q (\genblk1.pcpi_mul_rs2 [3]));
  DFFHQX1 \genblk1.pcpi_mul_rs2_reg[4] (.CK (clk), .D (n_1690), .Q
       (\genblk1.pcpi_mul_rs2 [4]));
  MDFFHQX4 \genblk1.pcpi_mul_rs2_reg[5] (.CK (clk), .D0
       (\reg_op2[5]_9674 ), .D1 (\genblk1.pcpi_mul_rs2 [5]), .S0
       (n_672), .Q (\genblk1.pcpi_mul_rs2 [5]));
  DFFHQX1 \genblk1.pcpi_mul_rs2_reg[6] (.CK (clk), .D (n_1680), .Q
       (\genblk1.pcpi_mul_rs2 [6]));
  MDFFHQX4 \genblk1.pcpi_mul_rs2_reg[7] (.CK (clk), .D0
       (\reg_op2[7]_9676 ), .D1 (\genblk1.pcpi_mul_rs2 [7]), .S0
       (n_672), .Q (\genblk1.pcpi_mul_rs2 [7]));
  DFFHQX1 \genblk1.pcpi_mul_rs2_reg[8] (.CK (clk), .D (n_1671), .Q
       (\genblk1.pcpi_mul_rs2 [8]));
  MDFFHQX4 \genblk1.pcpi_mul_rs2_reg[9] (.CK (clk), .D0
       (\reg_op2[9]_9678 ), .D1 (\genblk1.pcpi_mul_rs2 [9]), .S0
       (n_672), .Q (\genblk1.pcpi_mul_rs2 [9]));
  DFFHQX1 \genblk1.pcpi_mul_rs2_reg[10] (.CK (clk), .D (n_1673), .Q
       (\genblk1.pcpi_mul_rs2 [10]));
  MDFFHQX4 \genblk1.pcpi_mul_rs2_reg[11] (.CK (clk), .D0
       (\reg_op2[11]_9680 ), .D1 (\genblk1.pcpi_mul_rs2 [11]), .S0
       (n_672), .Q (\genblk1.pcpi_mul_rs2 [11]));
  DFFHQX1 \genblk1.pcpi_mul_rs2_reg[12] (.CK (clk), .D (n_1674), .Q
       (\genblk1.pcpi_mul_rs2 [12]));
  MDFFHQX4 \genblk1.pcpi_mul_rs2_reg[13] (.CK (clk), .D0
       (\reg_op2[13]_9682 ), .D1 (\genblk1.pcpi_mul_rs2 [13]), .S0
       (n_672), .Q (\genblk1.pcpi_mul_rs2 [13]));
  DFFHQX1 \genblk1.pcpi_mul_rs2_reg[14] (.CK (clk), .D (n_1689), .Q
       (\genblk1.pcpi_mul_rs2 [14]));
  MDFFHQX4 \genblk1.pcpi_mul_rs2_reg[15] (.CK (clk), .D0
       (\reg_op2[15]_9684 ), .D1 (\genblk1.pcpi_mul_rs2 [15]), .S0
       (n_672), .Q (\genblk1.pcpi_mul_rs2 [15]));
  DFFHQX1 \genblk1.pcpi_mul_rs2_reg[16] (.CK (clk), .D (n_1688), .Q
       (\genblk1.pcpi_mul_rs2 [16]));
  MDFFHQX4 \genblk1.pcpi_mul_rs2_reg[17] (.CK (clk), .D0
       (\reg_op2[17]_9686 ), .D1 (\genblk1.pcpi_mul_rs2 [17]), .S0
       (n_672), .Q (\genblk1.pcpi_mul_rs2 [17]));
  DFFHQX1 \genblk1.pcpi_mul_rs2_reg[18] (.CK (clk), .D (n_1687), .Q
       (\genblk1.pcpi_mul_rs2 [18]));
  MDFFHQX4 \genblk1.pcpi_mul_rs2_reg[19] (.CK (clk), .D0
       (\reg_op2[19]_9688 ), .D1 (\genblk1.pcpi_mul_rs2 [19]), .S0
       (n_672), .Q (\genblk1.pcpi_mul_rs2 [19]));
  DFFHQX1 \genblk1.pcpi_mul_rs2_reg[20] (.CK (clk), .D (n_1686), .Q
       (\genblk1.pcpi_mul_rs2 [20]));
  MDFFHQX4 \genblk1.pcpi_mul_rs2_reg[21] (.CK (clk), .D0
       (\reg_op2[21]_9690 ), .D1 (\genblk1.pcpi_mul_rs2 [21]), .S0
       (n_672), .Q (\genblk1.pcpi_mul_rs2 [21]));
  DFFHQX1 \genblk1.pcpi_mul_rs2_reg[22] (.CK (clk), .D (n_1685), .Q
       (\genblk1.pcpi_mul_rs2 [22]));
  MDFFHQX4 \genblk1.pcpi_mul_rs2_reg[23] (.CK (clk), .D0
       (\reg_op2[23]_9692 ), .D1 (\genblk1.pcpi_mul_rs2 [23]), .S0
       (n_672), .Q (\genblk1.pcpi_mul_rs2 [23]));
  DFFHQX1 \genblk1.pcpi_mul_rs2_reg[24] (.CK (clk), .D (n_1684), .Q
       (\genblk1.pcpi_mul_rs2 [24]));
  MDFFHQX4 \genblk1.pcpi_mul_rs2_reg[25] (.CK (clk), .D0
       (\reg_op2[25]_9694 ), .D1 (\genblk1.pcpi_mul_rs2 [25]), .S0
       (n_672), .Q (\genblk1.pcpi_mul_rs2 [25]));
  DFFHQX1 \genblk1.pcpi_mul_rs2_reg[26] (.CK (clk), .D (n_1683), .Q
       (\genblk1.pcpi_mul_rs2 [26]));
  MDFFHQX4 \genblk1.pcpi_mul_rs2_reg[27] (.CK (clk), .D0
       (\reg_op2[27]_9696 ), .D1 (\genblk1.pcpi_mul_rs2 [27]), .S0
       (n_672), .Q (\genblk1.pcpi_mul_rs2 [27]));
  DFFHQX1 \genblk1.pcpi_mul_rs2_reg[28] (.CK (clk), .D (n_1682), .Q
       (\genblk1.pcpi_mul_rs2 [28]));
  MDFFHQX4 \genblk1.pcpi_mul_rs2_reg[29] (.CK (clk), .D0
       (\reg_op2[29]_9698 ), .D1 (\genblk1.pcpi_mul_rs2 [29]), .S0
       (n_672), .Q (\genblk1.pcpi_mul_rs2 [29]));
  DFFHQX1 \genblk1.pcpi_mul_rs2_reg[30] (.CK (clk), .D (n_1681), .Q
       (\genblk1.pcpi_mul_rs2 [30]));
  MDFFHQX4 \genblk1.pcpi_mul_rs2_reg[31] (.CK (clk), .D0
       (\reg_op2[31]_9700 ), .D1 (\genblk1.pcpi_mul_rs2 [31]), .S0
       (n_672), .Q (\genblk1.pcpi_mul_rs2 [31]));
  DFFHQX1 \genblk2.pcpi_div_dividend_reg[0] (.CK (clk), .D (n_5497), .Q
       (\genblk2.pcpi_div_dividend [0]));
  DFFHQX1 \genblk2.pcpi_div_dividend_reg[1] (.CK (clk), .D (n_5496), .Q
       (\genblk2.pcpi_div_dividend [1]));
  DFFHQX1 \genblk2.pcpi_div_dividend_reg[2] (.CK (clk), .D (n_5495), .Q
       (\genblk2.pcpi_div_dividend [2]));
  DFFHQX1 \genblk2.pcpi_div_dividend_reg[3] (.CK (clk), .D (n_5494), .Q
       (\genblk2.pcpi_div_dividend [3]));
  DFFHQX1 \genblk2.pcpi_div_dividend_reg[4] (.CK (clk), .D (n_5492), .Q
       (\genblk2.pcpi_div_dividend [4]));
  DFFHQX1 \genblk2.pcpi_div_dividend_reg[5] (.CK (clk), .D (n_5493), .Q
       (\genblk2.pcpi_div_dividend [5]));
  DFFHQX1 \genblk2.pcpi_div_dividend_reg[6] (.CK (clk), .D (n_5491), .Q
       (\genblk2.pcpi_div_dividend [6]));
  DFFHQX1 \genblk2.pcpi_div_dividend_reg[7] (.CK (clk), .D (n_5490), .Q
       (\genblk2.pcpi_div_dividend [7]));
  DFFHQX1 \genblk2.pcpi_div_dividend_reg[8] (.CK (clk), .D (n_5489), .Q
       (\genblk2.pcpi_div_dividend [8]));
  DFFHQX1 \genblk2.pcpi_div_dividend_reg[9] (.CK (clk), .D (n_5487), .Q
       (\genblk2.pcpi_div_dividend [9]));
  DFFHQX1 \genblk2.pcpi_div_dividend_reg[10] (.CK (clk), .D (n_5488),
       .Q (\genblk2.pcpi_div_dividend [10]));
  DFFHQX1 \genblk2.pcpi_div_dividend_reg[11] (.CK (clk), .D (n_5486),
       .Q (\genblk2.pcpi_div_dividend [11]));
  DFFHQX1 \genblk2.pcpi_div_dividend_reg[12] (.CK (clk), .D (n_5485),
       .Q (\genblk2.pcpi_div_dividend [12]));
  DFFHQX1 \genblk2.pcpi_div_dividend_reg[13] (.CK (clk), .D (n_5484),
       .Q (\genblk2.pcpi_div_dividend [13]));
  DFFHQX1 \genblk2.pcpi_div_dividend_reg[14] (.CK (clk), .D (n_5498),
       .Q (\genblk2.pcpi_div_dividend [14]));
  DFFHQX1 \genblk2.pcpi_div_dividend_reg[15] (.CK (clk), .D (n_5482),
       .Q (\genblk2.pcpi_div_dividend [15]));
  DFFHQX1 \genblk2.pcpi_div_dividend_reg[16] (.CK (clk), .D (n_5481),
       .Q (\genblk2.pcpi_div_dividend [16]));
  DFFHQX1 \genblk2.pcpi_div_dividend_reg[17] (.CK (clk), .D (n_5480),
       .Q (\genblk2.pcpi_div_dividend [17]));
  DFFHQX1 \genblk2.pcpi_div_dividend_reg[18] (.CK (clk), .D (n_5479),
       .Q (\genblk2.pcpi_div_dividend [18]));
  DFFHQX1 \genblk2.pcpi_div_dividend_reg[19] (.CK (clk), .D (n_5478),
       .Q (\genblk2.pcpi_div_dividend [19]));
  DFFHQX1 \genblk2.pcpi_div_dividend_reg[20] (.CK (clk), .D (n_5476),
       .Q (\genblk2.pcpi_div_dividend [20]));
  DFFHQX1 \genblk2.pcpi_div_dividend_reg[21] (.CK (clk), .D (n_5474),
       .Q (\genblk2.pcpi_div_dividend [21]));
  DFFHQX1 \genblk2.pcpi_div_dividend_reg[22] (.CK (clk), .D (n_5477),
       .Q (\genblk2.pcpi_div_dividend [22]));
  DFFHQX1 \genblk2.pcpi_div_dividend_reg[23] (.CK (clk), .D (n_5475),
       .Q (\genblk2.pcpi_div_dividend [23]));
  DFFHQX1 \genblk2.pcpi_div_dividend_reg[24] (.CK (clk), .D (n_5473),
       .Q (\genblk2.pcpi_div_dividend [24]));
  DFFHQX1 \genblk2.pcpi_div_dividend_reg[25] (.CK (clk), .D (n_5472),
       .Q (\genblk2.pcpi_div_dividend [25]));
  DFFHQX1 \genblk2.pcpi_div_dividend_reg[26] (.CK (clk), .D (n_5471),
       .Q (\genblk2.pcpi_div_dividend [26]));
  DFFHQX1 \genblk2.pcpi_div_dividend_reg[27] (.CK (clk), .D (n_5470),
       .Q (\genblk2.pcpi_div_dividend [27]));
  DFFHQX1 \genblk2.pcpi_div_dividend_reg[28] (.CK (clk), .D (n_5469),
       .Q (\genblk2.pcpi_div_dividend [28]));
  DFFHQX1 \genblk2.pcpi_div_dividend_reg[29] (.CK (clk), .D (n_5468),
       .Q (\genblk2.pcpi_div_dividend [29]));
  DFFHQX1 \genblk2.pcpi_div_dividend_reg[30] (.CK (clk), .D (n_5467),
       .Q (\genblk2.pcpi_div_dividend [30]));
  DFFHQX1 \genblk2.pcpi_div_dividend_reg[31] (.CK (clk), .D (n_5466),
       .Q (\genblk2.pcpi_div_dividend [31]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[0] (.CK (clk), .D (n_5365), .Q
       (\genblk2.pcpi_div_divisor [0]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[1] (.CK (clk), .D (n_5364), .Q
       (\genblk2.pcpi_div_divisor [1]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[2] (.CK (clk), .D (n_5363), .Q
       (\genblk2.pcpi_div_divisor [2]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[3] (.CK (clk), .D (n_5362), .Q
       (\genblk2.pcpi_div_divisor [3]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[4] (.CK (clk), .D (n_5361), .Q
       (\genblk2.pcpi_div_divisor [4]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[5] (.CK (clk), .D (n_5360), .Q
       (\genblk2.pcpi_div_divisor [5]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[6] (.CK (clk), .D (n_5359), .Q
       (\genblk2.pcpi_div_divisor [6]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[7] (.CK (clk), .D (n_5358), .Q
       (\genblk2.pcpi_div_divisor [7]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[8] (.CK (clk), .D (n_5357), .Q
       (\genblk2.pcpi_div_divisor [8]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[9] (.CK (clk), .D (n_5356), .Q
       (\genblk2.pcpi_div_divisor [9]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[10] (.CK (clk), .D (n_5355), .Q
       (\genblk2.pcpi_div_divisor [10]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[11] (.CK (clk), .D (n_5354), .Q
       (\genblk2.pcpi_div_divisor [11]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[12] (.CK (clk), .D (n_5353), .Q
       (\genblk2.pcpi_div_divisor [12]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[13] (.CK (clk), .D (n_5352), .Q
       (\genblk2.pcpi_div_divisor [13]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[14] (.CK (clk), .D (n_5351), .Q
       (\genblk2.pcpi_div_divisor [14]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[15] (.CK (clk), .D (n_5349), .Q
       (\genblk2.pcpi_div_divisor [15]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[16] (.CK (clk), .D (n_5350), .Q
       (\genblk2.pcpi_div_divisor [16]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[17] (.CK (clk), .D (n_5348), .Q
       (\genblk2.pcpi_div_divisor [17]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[18] (.CK (clk), .D (n_5347), .Q
       (\genblk2.pcpi_div_divisor [18]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[19] (.CK (clk), .D (n_5346), .Q
       (\genblk2.pcpi_div_divisor [19]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[20] (.CK (clk), .D (n_5345), .Q
       (\genblk2.pcpi_div_divisor [20]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[21] (.CK (clk), .D (n_5344), .Q
       (\genblk2.pcpi_div_divisor [21]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[22] (.CK (clk), .D (n_5366), .Q
       (\genblk2.pcpi_div_divisor [22]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[23] (.CK (clk), .D (n_5342), .Q
       (\genblk2.pcpi_div_divisor [23]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[24] (.CK (clk), .D (n_5341), .Q
       (\genblk2.pcpi_div_divisor [24]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[25] (.CK (clk), .D (n_5340), .Q
       (\genblk2.pcpi_div_divisor [25]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[26] (.CK (clk), .D (n_5339), .Q
       (\genblk2.pcpi_div_divisor [26]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[27] (.CK (clk), .D (n_5338), .Q
       (\genblk2.pcpi_div_divisor [27]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[28] (.CK (clk), .D (n_5337), .Q
       (\genblk2.pcpi_div_divisor [28]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[29] (.CK (clk), .D (n_5336), .Q
       (\genblk2.pcpi_div_divisor [29]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[30] (.CK (clk), .D (n_5335), .Q
       (\genblk2.pcpi_div_divisor [30]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[31] (.CK (clk), .D (n_5399), .Q
       (\genblk2.pcpi_div_divisor [31]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[32] (.CK (clk), .D (n_5425), .Q
       (\genblk2.pcpi_div_divisor [32]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[33] (.CK (clk), .D (n_5424), .Q
       (\genblk2.pcpi_div_divisor [33]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[34] (.CK (clk), .D (n_5423), .Q
       (\genblk2.pcpi_div_divisor [34]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[35] (.CK (clk), .D (n_5422), .Q
       (\genblk2.pcpi_div_divisor [35]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[36] (.CK (clk), .D (n_5421), .Q
       (\genblk2.pcpi_div_divisor [36]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[37] (.CK (clk), .D (n_5420), .Q
       (\genblk2.pcpi_div_divisor [37]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[38] (.CK (clk), .D (n_5419), .Q
       (\genblk2.pcpi_div_divisor [38]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[39] (.CK (clk), .D (n_5417), .Q
       (\genblk2.pcpi_div_divisor [39]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[40] (.CK (clk), .D (n_5418), .Q
       (\genblk2.pcpi_div_divisor [40]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[41] (.CK (clk), .D (n_5416), .Q
       (\genblk2.pcpi_div_divisor [41]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[42] (.CK (clk), .D (n_5415), .Q
       (\genblk2.pcpi_div_divisor [42]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[43] (.CK (clk), .D (n_5414), .Q
       (\genblk2.pcpi_div_divisor [43]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[44] (.CK (clk), .D (n_5413), .Q
       (\genblk2.pcpi_div_divisor [44]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[45] (.CK (clk), .D (n_5412), .Q
       (\genblk2.pcpi_div_divisor [45]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[46] (.CK (clk), .D (n_5411), .Q
       (\genblk2.pcpi_div_divisor [46]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[47] (.CK (clk), .D (n_5410), .Q
       (\genblk2.pcpi_div_divisor [47]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[48] (.CK (clk), .D (n_5409), .Q
       (\genblk2.pcpi_div_divisor [48]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[49] (.CK (clk), .D (n_5408), .Q
       (\genblk2.pcpi_div_divisor [49]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[50] (.CK (clk), .D (n_5400), .Q
       (\genblk2.pcpi_div_divisor [50]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[51] (.CK (clk), .D (n_5407), .Q
       (\genblk2.pcpi_div_divisor [51]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[52] (.CK (clk), .D (n_5429), .Q
       (\genblk2.pcpi_div_divisor [52]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[53] (.CK (clk), .D (n_5428), .Q
       (\genblk2.pcpi_div_divisor [53]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[54] (.CK (clk), .D (n_5427), .Q
       (\genblk2.pcpi_div_divisor [54]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[55] (.CK (clk), .D (n_5406), .Q
       (\genblk2.pcpi_div_divisor [55]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[56] (.CK (clk), .D (n_5405), .Q
       (\genblk2.pcpi_div_divisor [56]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[57] (.CK (clk), .D (n_5404), .Q
       (\genblk2.pcpi_div_divisor [57]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[58] (.CK (clk), .D (n_5403), .Q
       (\genblk2.pcpi_div_divisor [58]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[59] (.CK (clk), .D (n_5402), .Q
       (\genblk2.pcpi_div_divisor [59]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[60] (.CK (clk), .D (n_5401), .Q
       (\genblk2.pcpi_div_divisor [60]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[61] (.CK (clk), .D (n_5426), .Q
       (\genblk2.pcpi_div_divisor [61]));
  DFFHQX1 \genblk2.pcpi_div_divisor_reg[62] (.CK (clk), .D (n_5398), .Q
       (\genblk2.pcpi_div_divisor [62]));
  DFFHQX1 \genblk2.pcpi_div_pcpi_ready_reg (.CK (clk), .D (n_5265), .Q
       (pcpi_div_wr));
  DFFHQX1 \genblk2.pcpi_div_quotient_msk_reg[0] (.CK (clk), .D
       (n_5302), .Q (\genblk2.pcpi_div_quotient_msk [0]));
  DFFHQX1 \genblk2.pcpi_div_quotient_msk_reg[1] (.CK (clk), .D
       (n_5301), .Q (\genblk2.pcpi_div_quotient_msk [1]));
  DFFHQX1 \genblk2.pcpi_div_quotient_msk_reg[2] (.CK (clk), .D
       (n_5300), .Q (\genblk2.pcpi_div_quotient_msk [2]));
  DFFHQX1 \genblk2.pcpi_div_quotient_msk_reg[3] (.CK (clk), .D
       (n_5299), .Q (\genblk2.pcpi_div_quotient_msk [3]));
  DFFHQX1 \genblk2.pcpi_div_quotient_msk_reg[4] (.CK (clk), .D
       (n_5298), .Q (\genblk2.pcpi_div_quotient_msk [4]));
  DFFHQX1 \genblk2.pcpi_div_quotient_msk_reg[5] (.CK (clk), .D
       (n_5291), .Q (\genblk2.pcpi_div_quotient_msk [5]));
  DFFHQX1 \genblk2.pcpi_div_quotient_msk_reg[6] (.CK (clk), .D
       (n_5295), .Q (\genblk2.pcpi_div_quotient_msk [6]));
  DFFHQX1 \genblk2.pcpi_div_quotient_msk_reg[7] (.CK (clk), .D
       (n_5297), .Q (\genblk2.pcpi_div_quotient_msk [7]));
  DFFHQX1 \genblk2.pcpi_div_quotient_msk_reg[8] (.CK (clk), .D
       (n_5296), .Q (\genblk2.pcpi_div_quotient_msk [8]));
  DFFHQX1 \genblk2.pcpi_div_quotient_msk_reg[9] (.CK (clk), .D
       (n_5294), .Q (\genblk2.pcpi_div_quotient_msk [9]));
  DFFHQX1 \genblk2.pcpi_div_quotient_msk_reg[10] (.CK (clk), .D
       (n_5293), .Q (\genblk2.pcpi_div_quotient_msk [10]));
  DFFHQX1 \genblk2.pcpi_div_quotient_msk_reg[11] (.CK (clk), .D
       (n_5292), .Q (\genblk2.pcpi_div_quotient_msk [11]));
  DFFHQX1 \genblk2.pcpi_div_quotient_msk_reg[12] (.CK (clk), .D
       (n_5290), .Q (\genblk2.pcpi_div_quotient_msk [12]));
  DFFHQX1 \genblk2.pcpi_div_quotient_msk_reg[13] (.CK (clk), .D
       (n_5289), .Q (\genblk2.pcpi_div_quotient_msk [13]));
  DFFHQX1 \genblk2.pcpi_div_quotient_msk_reg[14] (.CK (clk), .D
       (n_5288), .Q (\genblk2.pcpi_div_quotient_msk [14]));
  DFFHQX1 \genblk2.pcpi_div_quotient_msk_reg[15] (.CK (clk), .D
       (n_5287), .Q (\genblk2.pcpi_div_quotient_msk [15]));
  DFFHQX1 \genblk2.pcpi_div_quotient_msk_reg[16] (.CK (clk), .D
       (n_5286), .Q (\genblk2.pcpi_div_quotient_msk [16]));
  DFFHQX1 \genblk2.pcpi_div_quotient_msk_reg[17] (.CK (clk), .D
       (n_5285), .Q (\genblk2.pcpi_div_quotient_msk [17]));
  DFFHQX1 \genblk2.pcpi_div_quotient_msk_reg[18] (.CK (clk), .D
       (n_5284), .Q (\genblk2.pcpi_div_quotient_msk [18]));
  DFFHQX1 \genblk2.pcpi_div_quotient_msk_reg[19] (.CK (clk), .D
       (n_5283), .Q (\genblk2.pcpi_div_quotient_msk [19]));
  DFFHQX1 \genblk2.pcpi_div_quotient_msk_reg[20] (.CK (clk), .D
       (n_5282), .Q (\genblk2.pcpi_div_quotient_msk [20]));
  DFFHQX1 \genblk2.pcpi_div_quotient_msk_reg[21] (.CK (clk), .D
       (n_5279), .Q (\genblk2.pcpi_div_quotient_msk [21]));
  DFFHQX1 \genblk2.pcpi_div_quotient_msk_reg[22] (.CK (clk), .D
       (n_5281), .Q (\genblk2.pcpi_div_quotient_msk [22]));
  DFFHQX1 \genblk2.pcpi_div_quotient_msk_reg[23] (.CK (clk), .D
       (n_5280), .Q (\genblk2.pcpi_div_quotient_msk [23]));
  DFFHQX1 \genblk2.pcpi_div_quotient_msk_reg[24] (.CK (clk), .D
       (n_5278), .Q (\genblk2.pcpi_div_quotient_msk [24]));
  DFFHQX1 \genblk2.pcpi_div_quotient_msk_reg[25] (.CK (clk), .D
       (n_5277), .Q (\genblk2.pcpi_div_quotient_msk [25]));
  DFFHQX1 \genblk2.pcpi_div_quotient_msk_reg[26] (.CK (clk), .D
       (n_5276), .Q (\genblk2.pcpi_div_quotient_msk [26]));
  DFFHQX1 \genblk2.pcpi_div_quotient_msk_reg[27] (.CK (clk), .D
       (n_5275), .Q (\genblk2.pcpi_div_quotient_msk [27]));
  DFFHQX1 \genblk2.pcpi_div_quotient_msk_reg[28] (.CK (clk), .D
       (n_5274), .Q (\genblk2.pcpi_div_quotient_msk [28]));
  DFFHQX1 \genblk2.pcpi_div_quotient_msk_reg[29] (.CK (clk), .D
       (n_5273), .Q (\genblk2.pcpi_div_quotient_msk [29]));
  DFFHQX1 \genblk2.pcpi_div_quotient_msk_reg[30] (.CK (clk), .D
       (n_5272), .Q (\genblk2.pcpi_div_quotient_msk [30]));
  DFFHQX1 \genblk2.pcpi_div_quotient_msk_reg[31] (.CK (clk), .D
       (n_5343), .Q (\genblk2.pcpi_div_quotient_msk [31]));
  DFFHQX1 \genblk2.pcpi_div_quotient_reg[0] (.CK (clk), .D (n_11768),
       .Q (\genblk2.pcpi_div_quotient [0]));
  DFFHQX1 \genblk2.pcpi_div_quotient_reg[1] (.CK (clk), .D (n_11769),
       .Q (\genblk2.pcpi_div_quotient [1]));
  DFFHQX1 \genblk2.pcpi_div_quotient_reg[2] (.CK (clk), .D (n_11770),
       .Q (\genblk2.pcpi_div_quotient [2]));
  DFFHQX1 \genblk2.pcpi_div_quotient_reg[3] (.CK (clk), .D (n_11771),
       .Q (\genblk2.pcpi_div_quotient [3]));
  DFFHQX1 \genblk2.pcpi_div_quotient_reg[4] (.CK (clk), .D (n_11772),
       .Q (\genblk2.pcpi_div_quotient [4]));
  DFFHQX1 \genblk2.pcpi_div_quotient_reg[5] (.CK (clk), .D (n_11773),
       .Q (\genblk2.pcpi_div_quotient [5]));
  DFFHQX1 \genblk2.pcpi_div_quotient_reg[6] (.CK (clk), .D (n_11775),
       .Q (\genblk2.pcpi_div_quotient [6]));
  DFFHQX1 \genblk2.pcpi_div_quotient_reg[7] (.CK (clk), .D (n_11774),
       .Q (\genblk2.pcpi_div_quotient [7]));
  DFFHQX1 \genblk2.pcpi_div_quotient_reg[8] (.CK (clk), .D (n_11776),
       .Q (\genblk2.pcpi_div_quotient [8]));
  DFFHQX1 \genblk2.pcpi_div_quotient_reg[9] (.CK (clk), .D (n_11777),
       .Q (\genblk2.pcpi_div_quotient [9]));
  DFFHQX1 \genblk2.pcpi_div_quotient_reg[10] (.CK (clk), .D (n_11778),
       .Q (\genblk2.pcpi_div_quotient [10]));
  DFFHQX1 \genblk2.pcpi_div_quotient_reg[11] (.CK (clk), .D (n_11779),
       .Q (\genblk2.pcpi_div_quotient [11]));
  DFFHQX1 \genblk2.pcpi_div_quotient_reg[12] (.CK (clk), .D (n_11780),
       .Q (\genblk2.pcpi_div_quotient [12]));
  DFFHQX1 \genblk2.pcpi_div_quotient_reg[13] (.CK (clk), .D (n_11781),
       .Q (\genblk2.pcpi_div_quotient [13]));
  DFFHQX1 \genblk2.pcpi_div_quotient_reg[14] (.CK (clk), .D (n_11782),
       .Q (\genblk2.pcpi_div_quotient [14]));
  DFFHQX1 \genblk2.pcpi_div_quotient_reg[15] (.CK (clk), .D (n_11783),
       .Q (\genblk2.pcpi_div_quotient [15]));
  DFFHQX1 \genblk2.pcpi_div_quotient_reg[16] (.CK (clk), .D (n_11784),
       .Q (\genblk2.pcpi_div_quotient [16]));
  DFFHQX1 \genblk2.pcpi_div_quotient_reg[17] (.CK (clk), .D (n_11785),
       .Q (\genblk2.pcpi_div_quotient [17]));
  DFFHQX1 \genblk2.pcpi_div_quotient_reg[18] (.CK (clk), .D (n_11786),
       .Q (\genblk2.pcpi_div_quotient [18]));
  DFFHQX1 \genblk2.pcpi_div_quotient_reg[19] (.CK (clk), .D (n_11787),
       .Q (\genblk2.pcpi_div_quotient [19]));
  DFFHQX1 \genblk2.pcpi_div_quotient_reg[20] (.CK (clk), .D (n_11788),
       .Q (\genblk2.pcpi_div_quotient [20]));
  DFFHQX1 \genblk2.pcpi_div_quotient_reg[21] (.CK (clk), .D (n_11791),
       .Q (\genblk2.pcpi_div_quotient [21]));
  DFFHQX1 \genblk2.pcpi_div_quotient_reg[22] (.CK (clk), .D (n_11789),
       .Q (\genblk2.pcpi_div_quotient [22]));
  DFFHQX1 \genblk2.pcpi_div_quotient_reg[23] (.CK (clk), .D (n_11790),
       .Q (\genblk2.pcpi_div_quotient [23]));
  DFFHQX1 \genblk2.pcpi_div_quotient_reg[24] (.CK (clk), .D (n_11792),
       .Q (\genblk2.pcpi_div_quotient [24]));
  DFFHQX1 \genblk2.pcpi_div_quotient_reg[25] (.CK (clk), .D (n_11793),
       .Q (\genblk2.pcpi_div_quotient [25]));
  DFFHQX1 \genblk2.pcpi_div_quotient_reg[26] (.CK (clk), .D (n_11794),
       .Q (\genblk2.pcpi_div_quotient [26]));
  DFFHQX1 \genblk2.pcpi_div_quotient_reg[27] (.CK (clk), .D (n_11795),
       .Q (\genblk2.pcpi_div_quotient [27]));
  DFFHQX1 \genblk2.pcpi_div_quotient_reg[28] (.CK (clk), .D (n_11796),
       .Q (\genblk2.pcpi_div_quotient [28]));
  DFFHQX1 \genblk2.pcpi_div_quotient_reg[29] (.CK (clk), .D (n_11797),
       .Q (\genblk2.pcpi_div_quotient [29]));
  DFFHQX1 \genblk2.pcpi_div_quotient_reg[30] (.CK (clk), .D (n_11798),
       .Q (\genblk2.pcpi_div_quotient [30]));
  DFFHQX1 \genblk2.pcpi_div_quotient_reg[31] (.CK (clk), .D (n_11767),
       .Q (\genblk2.pcpi_div_quotient [31]));
  DFFHQX1 \genblk2.pcpi_div_running_reg (.CK (clk), .D (n_5268), .Q
       (\genblk2.pcpi_div_running ));
  DFFHQX1 instr_add_reg(.CK (clk), .D (n_2973), .Q (instr_add));
  DFFHQX1 instr_addi_reg(.CK (clk), .D (n_2282), .Q (instr_addi));
  DFFHQX1 instr_and_reg(.CK (clk), .D (n_2972), .Q (instr_and));
  DFFHQX1 instr_andi_reg(.CK (clk), .D (n_2283), .Q (instr_andi));
  DFFHQX1 instr_auipc_reg(.CK (clk), .D (n_3016), .Q (instr_auipc));
  DFFHQX1 instr_beq_reg(.CK (clk), .D (n_2284), .Q (instr_beq));
  DFFHQX1 instr_bge_reg(.CK (clk), .D (n_2285), .Q (instr_bge));
  DFFHQX1 instr_bgeu_reg(.CK (clk), .D (n_2286), .Q (instr_bgeu));
  DFFHQX1 instr_blt_reg(.CK (clk), .D (n_2287), .Q (instr_blt));
  DFFHQX1 instr_bltu_reg(.CK (clk), .D (n_2288), .Q (instr_bltu));
  DFFHQX1 instr_bne_reg(.CK (clk), .D (n_2289), .Q (instr_bne));
  DFFHQX1 instr_ecall_ebreak_reg(.CK (clk), .D (n_5084), .Q
       (instr_ecall_ebreak));
  DFFHQX1 instr_jalr_reg(.CK (clk), .D (n_4790), .Q (instr_jalr));
  DFFHQX1 instr_lb_reg(.CK (clk), .D (n_1992), .Q (instr_lb));
  DFFHQX1 instr_lbu_reg(.CK (clk), .D (n_1984), .Q (instr_lbu));
  DFFHQX1 instr_lh_reg(.CK (clk), .D (n_1996), .Q (instr_lh));
  DFFHQX1 instr_lhu_reg(.CK (clk), .D (n_1990), .Q (instr_lhu));
  DFFHQX1 instr_lui_reg(.CK (clk), .D (n_4097), .Q (instr_lui));
  DFFHQX1 instr_lw_reg(.CK (clk), .D (n_1983), .Q (instr_lw));
  DFFHQX1 instr_or_reg(.CK (clk), .D (n_2970), .Q (instr_or));
  DFFHQX1 instr_ori_reg(.CK (clk), .D (n_2291), .Q (instr_ori));
  DFFQX2 instr_rdcycle_reg(.CK (clk), .D (n_4979), .Q (instr_rdcycle));
  DFFQX2 instr_rdcycleh_reg(.CK (clk), .D (n_5012), .Q
       (instr_rdcycleh));
  DFFQX2 instr_rdinstr_reg(.CK (clk), .D (n_5082), .Q (instr_rdinstr));
  DFFHQX1 instr_sb_reg(.CK (clk), .D (n_1991), .Q (instr_sb));
  DFFHQX1 instr_sh_reg(.CK (clk), .D (n_1995), .Q (instr_sh));
  DFFHQX1 instr_sll_reg(.CK (clk), .D (n_2969), .Q (instr_sll));
  DFFHQX1 instr_slli_reg(.CK (clk), .D (n_2570), .Q (instr_slli));
  DFFHQX1 instr_slt_reg(.CK (clk), .D (n_2968), .Q (instr_slt));
  DFFHQX1 instr_slti_reg(.CK (clk), .D (n_2292), .Q (instr_slti));
  DFFHQX1 instr_sltiu_reg(.CK (clk), .D (n_2312), .Q (instr_sltiu));
  DFFHQX1 instr_sltu_reg(.CK (clk), .D (n_3047), .Q (instr_sltu));
  DFFHQX1 instr_sra_reg(.CK (clk), .D (n_2967), .Q (instr_sra));
  DFFHQX1 instr_srai_reg(.CK (clk), .D (n_2560), .Q (instr_srai));
  DFFHQX1 instr_srl_reg(.CK (clk), .D (n_2966), .Q (instr_srl));
  DFFHQX1 instr_srli_reg(.CK (clk), .D (n_2573), .Q (instr_srli));
  DFFHQX1 instr_sw_reg(.CK (clk), .D (n_1980), .Q (instr_sw));
  DFFHQX1 instr_xor_reg(.CK (clk), .D (n_2964), .Q (instr_xor));
  DFFHQX1 instr_xori_reg(.CK (clk), .D (n_2294), .Q (instr_xori));
  DFFHQX1 is_alu_reg_reg_reg(.CK (clk), .D (n_3429), .Q
       (is_alu_reg_reg));
  DFFHQX1 is_beq_bne_blt_bge_bltu_bgeu_reg(.CK (clk), .D (n_3039), .Q
       (is_beq_bne_blt_bge_bltu_bgeu));
  DFFHQX1 is_jalr_addi_slti_sltiu_xori_ori_andi_reg(.CK (clk), .D
       (n_2363), .Q (is_jalr_addi_slti_sltiu_xori_ori_andi));
  DFFHQX1 is_lb_lh_lw_lbu_lhu_reg(.CK (clk), .D (n_3424), .Q
       (is_lb_lh_lw_lbu_lhu));
  DFFHQX1 is_sb_sh_sw_reg(.CK (clk), .D (n_3076), .Q (is_sb_sh_sw));
  DFFHQX1 is_sll_srl_sra_reg(.CK (clk), .D (n_3012), .Q
       (is_sll_srl_sra));
  DFFQX2 latched_branch_reg(.CK (clk), .D (n_5526), .Q
       (latched_branch));
  DFFHQX1 latched_compr_reg(.CK (clk), .D (n_1482), .Q (latched_compr));
  DFFHQX1 latched_is_lb_reg(.CK (clk), .D (n_2431), .Q (latched_is_lb));
  DFFHQX1 latched_is_lh_reg(.CK (clk), .D (n_2428), .Q (latched_is_lh));
  DFFHQX1 latched_is_lu_reg(.CK (clk), .D (n_2429), .Q (latched_is_lu));
  DFFHQX1 \latched_rd_reg[0] (.CK (clk), .D (n_1743), .Q
       (latched_rd[0]));
  DFFQX2 latched_stalu_reg(.CK (clk), .D (n_2161), .Q (latched_stalu));
  DFFHQX1 latched_store_reg(.CK (clk), .D (n_5527), .Q (latched_store));
  DFFHQX1 \mem_16bit_buffer_reg[0] (.CK (clk), .D (n_2551), .Q
       (mem_16bit_buffer[0]));
  DFFHQX1 \mem_16bit_buffer_reg[1] (.CK (clk), .D (n_2550), .Q
       (mem_16bit_buffer[1]));
  DFFHQX1 \mem_16bit_buffer_reg[2] (.CK (clk), .D (n_2549), .Q
       (mem_16bit_buffer[2]));
  DFFHQX1 \mem_16bit_buffer_reg[3] (.CK (clk), .D (n_2548), .Q
       (mem_16bit_buffer[3]));
  DFFHQX1 \mem_16bit_buffer_reg[4] (.CK (clk), .D (n_2547), .Q
       (mem_16bit_buffer[4]));
  DFFHQX1 \mem_16bit_buffer_reg[5] (.CK (clk), .D (n_2546), .Q
       (mem_16bit_buffer[5]));
  DFFHQX1 \mem_16bit_buffer_reg[6] (.CK (clk), .D (n_2545), .Q
       (mem_16bit_buffer[6]));
  DFFHQX1 \mem_16bit_buffer_reg[7] (.CK (clk), .D (n_2544), .Q
       (mem_16bit_buffer[7]));
  DFFHQX1 \mem_16bit_buffer_reg[8] (.CK (clk), .D (n_2543), .Q
       (mem_16bit_buffer[8]));
  DFFHQX1 \mem_16bit_buffer_reg[9] (.CK (clk), .D (n_2542), .Q
       (mem_16bit_buffer[9]));
  DFFHQX1 \mem_16bit_buffer_reg[10] (.CK (clk), .D (n_2541), .Q
       (mem_16bit_buffer[10]));
  DFFHQX1 \mem_16bit_buffer_reg[11] (.CK (clk), .D (n_2540), .Q
       (mem_16bit_buffer[11]));
  DFFHQX1 \mem_16bit_buffer_reg[12] (.CK (clk), .D (n_2539), .Q
       (mem_16bit_buffer[12]));
  DFFHQX1 \mem_16bit_buffer_reg[13] (.CK (clk), .D (n_2538), .Q
       (mem_16bit_buffer[13]));
  DFFHQX1 \mem_16bit_buffer_reg[14] (.CK (clk), .D (n_2537), .Q
       (mem_16bit_buffer[14]));
  DFFHQX1 \mem_16bit_buffer_reg[15] (.CK (clk), .D (n_2536), .Q
       (mem_16bit_buffer[15]));
  DFFHQX1 \mem_addr_reg[2] (.CK (clk), .D (n_8829), .Q (n_5662));
  DFFHQX1 \mem_addr_reg[3] (.CK (clk), .D (n_9060), .Q (n_5663));
  DFFHQX1 \mem_addr_reg[4] (.CK (clk), .D (n_9039), .Q (n_5664));
  DFFHQX1 \mem_addr_reg[5] (.CK (clk), .D (n_9018), .Q (n_5665));
  DFFHQX1 \mem_addr_reg[6] (.CK (clk), .D (n_9354), .Q (n_5666));
  DFFHQX1 \mem_addr_reg[7] (.CK (clk), .D (n_8997), .Q (n_5667));
  DFFHQX1 \mem_addr_reg[8] (.CK (clk), .D (n_8955), .Q (n_5668));
  DFFHQX1 \mem_addr_reg[9] (.CK (clk), .D (n_8934), .Q (n_5669));
  DFFHQX1 \mem_addr_reg[10] (.CK (clk), .D (n_9438), .Q (n_5670));
  DFFHQX1 \mem_addr_reg[11] (.CK (clk), .D (n_8913), .Q (n_5671));
  DFFHQX1 \mem_addr_reg[12] (.CK (clk), .D (n_8871), .Q (n_5672));
  DFFHQX1 \mem_addr_reg[13] (.CK (clk), .D (n_8850), .Q (n_5673));
  DFFHQX1 \mem_addr_reg[14] (.CK (clk), .D (n_9417), .Q (n_5674));
  DFFHQX1 \mem_addr_reg[15] (.CK (clk), .D (n_8787), .Q (n_5675));
  DFFHQX1 \mem_addr_reg[16] (.CK (clk), .D (n_8766), .Q (n_5676));
  DFFHQX1 \mem_addr_reg[17] (.CK (clk), .D (n_8745), .Q (n_5677));
  DFFHQX1 \mem_addr_reg[18] (.CK (clk), .D (n_8556), .Q (n_5678));
  DFFHQX1 \mem_addr_reg[19] (.CK (clk), .D (n_8724), .Q (n_5679));
  DFFHQX1 \mem_addr_reg[20] (.CK (clk), .D (n_8703), .Q (n_5680));
  DFFHQX1 \mem_addr_reg[21] (.CK (clk), .D (n_8682), .Q (n_5681));
  DFFHQX1 \mem_addr_reg[22] (.CK (clk), .D (n_8661), .Q (n_5682));
  DFFHQX1 \mem_addr_reg[23] (.CK (clk), .D (n_8640), .Q (n_5683));
  DFFHQX1 \mem_addr_reg[24] (.CK (clk), .D (n_8619), .Q (n_5684));
  DFFHQX1 \mem_addr_reg[25] (.CK (clk), .D (n_8598), .Q (n_5685));
  DFFHQX1 \mem_addr_reg[26] (.CK (clk), .D (n_8577), .Q (n_5686));
  DFFHQX1 \mem_addr_reg[27] (.CK (clk), .D (n_8535), .Q (n_5687));
  DFFHQX1 \mem_addr_reg[28] (.CK (clk), .D (n_8514), .Q (n_5688));
  DFFHQX1 \mem_addr_reg[29] (.CK (clk), .D (n_8493), .Q (n_5689));
  DFFHQX1 \mem_addr_reg[30] (.CK (clk), .D (n_8808), .Q (n_5690));
  DFFHQX1 \mem_addr_reg[31] (.CK (clk), .D (n_9690), .Q (n_5691));
  DFFHQX1 mem_do_wdata_reg(.CK (clk), .D (n_2344), .Q (mem_do_wdata));
  DFFHQX1 mem_instr_reg(.CK (clk), .D (n_2104), .Q (n_5692));
  DFFHQX1 mem_la_firstword_reg_reg(.CK (clk), .D (n_1550), .Q
       (mem_la_firstword_reg));
  DFFHQX1 mem_la_secondword_reg(.CK (clk), .D (n_2125), .Q
       (mem_la_secondword));
  DFFHQX1 \mem_rdata_q_reg[0] (.CK (clk), .D (n_994), .Q
       (mem_rdata_q[0]));
  DFFHQX1 \mem_rdata_q_reg[1] (.CK (clk), .D (n_1027), .Q
       (mem_rdata_q[1]));
  DFFHQX1 \mem_rdata_q_reg[2] (.CK (clk), .D (n_2343), .Q
       (mem_rdata_q[2]));
  DFFHQX1 \mem_rdata_q_reg[3] (.CK (clk), .D (n_11799), .Q
       (mem_rdata_q[3]));
  DFFHQX1 \mem_rdata_q_reg[10] (.CK (clk), .D (n_3260), .Q
       (mem_rdata_q[10]));
  DFFHQX1 \mem_rdata_q_reg[11] (.CK (clk), .D (n_3259), .Q
       (mem_rdata_q[11]));
  DFFHQX1 \mem_rdata_q_reg[16] (.CK (clk), .D (n_4715), .Q
       (mem_rdata_q[16]));
  DFFHQX1 \mem_rdata_q_reg[17] (.CK (clk), .D (n_4773), .Q
       (mem_rdata_q[17]));
  DFFHQX1 \mem_rdata_q_reg[28] (.CK (clk), .D (n_5198), .Q
       (mem_rdata_q[28]));
  DFFHQX1 \mem_rdata_q_reg[29] (.CK (clk), .D (n_5168), .Q
       (mem_rdata_q[29]));
  DFFHQX1 \mem_state_reg[0] (.CK (clk), .D (n_3172), .Q (mem_state[0]));
  DFFHQX1 mem_valid_reg(.CK (clk), .D (n_2947), .Q (mem_valid_9465));
  DFFHQX1 \mem_wdata_reg[0] (.CK (clk), .D (n_1661), .Q (n_5630));
  DFFHQX1 \mem_wdata_reg[1] (.CK (clk), .D (n_1660), .Q (n_5631));
  DFFHQX1 \mem_wdata_reg[2] (.CK (clk), .D (n_1659), .Q (n_5632));
  DFFHQX1 \mem_wdata_reg[3] (.CK (clk), .D (n_1658), .Q (n_5633));
  DFFHQX1 \mem_wdata_reg[4] (.CK (clk), .D (n_1657), .Q (n_5634));
  DFFHQX1 \mem_wdata_reg[5] (.CK (clk), .D (n_1656), .Q (n_5635));
  DFFHQX1 \mem_wdata_reg[6] (.CK (clk), .D (n_1655), .Q (n_5636));
  DFFHQX1 \mem_wdata_reg[7] (.CK (clk), .D (n_1654), .Q (n_5637));
  DFFHQX1 \mem_wdata_reg[8] (.CK (clk), .D (n_9669), .Q (n_5638));
  DFFHQX1 \mem_wdata_reg[9] (.CK (clk), .D (n_9648), .Q (n_5639));
  DFFHQX1 \mem_wdata_reg[10] (.CK (clk), .D (n_8892), .Q (n_5640));
  DFFHQX1 \mem_wdata_reg[11] (.CK (clk), .D (n_9627), .Q (n_5641));
  DFFHQX1 \mem_wdata_reg[12] (.CK (clk), .D (n_9606), .Q (n_5642));
  DFFHQX1 \mem_wdata_reg[13] (.CK (clk), .D (n_9585), .Q (n_5643));
  DFFHQX1 \mem_wdata_reg[14] (.CK (clk), .D (n_8976), .Q (n_5644));
  DFFHQX1 \mem_wdata_reg[15] (.CK (clk), .D (n_9564), .Q (n_5645));
  DFFHQX1 \mem_wdata_reg[16] (.CK (clk), .D (n_9165), .Q (n_5646));
  DFFHQX1 \mem_wdata_reg[17] (.CK (clk), .D (n_9543), .Q (n_5647));
  DFFHQX1 \mem_wdata_reg[18] (.CK (clk), .D (n_9228), .Q (n_5648));
  DFFHQX1 \mem_wdata_reg[19] (.CK (clk), .D (n_9501), .Q (n_5649));
  DFFHQX1 \mem_wdata_reg[20] (.CK (clk), .D (n_9207), .Q (n_5650));
  DFFHQX1 \mem_wdata_reg[21] (.CK (clk), .D (n_9522), .Q (n_5651));
  DFFHQX1 \mem_wdata_reg[22] (.CK (clk), .D (n_9249), .Q (n_5652));
  DFFHQX1 \mem_wdata_reg[23] (.CK (clk), .D (n_9186), .Q (n_5653));
  DFFHQX1 \mem_wdata_reg[24] (.CK (clk), .D (n_9291), .Q (n_5654));
  DFFHQX1 \mem_wdata_reg[25] (.CK (clk), .D (n_9480), .Q (n_5655));
  DFFHQX1 \mem_wdata_reg[26] (.CK (clk), .D (n_9333), .Q (n_5656));
  DFFHQX1 \mem_wdata_reg[27] (.CK (clk), .D (n_9312), .Q (n_5657));
  DFFHQX1 \mem_wdata_reg[28] (.CK (clk), .D (n_9459), .Q (n_5658));
  DFFHQX1 \mem_wdata_reg[29] (.CK (clk), .D (n_9270), .Q (n_5659));
  DFFHQX1 \mem_wdata_reg[30] (.CK (clk), .D (n_9375), .Q (n_5660));
  DFFHQX1 \mem_wdata_reg[31] (.CK (clk), .D (n_9396), .Q (n_5661));
  DFFHQX1 \mem_wordsize_reg[0] (.CK (clk), .D (n_2486), .Q
       (mem_wordsize[0]));
  DFFHQX1 \mem_wordsize_reg[1] (.CK (clk), .D (n_2487), .Q
       (mem_wordsize[1]));
  DFFHQX1 \mem_wstrb_reg[0] (.CK (clk), .D (n_9144), .Q (n_5626));
  DFFHQX1 \mem_wstrb_reg[1] (.CK (clk), .D (n_9123), .Q (n_5627));
  DFFHQX1 \mem_wstrb_reg[2] (.CK (clk), .D (n_9102), .Q (n_5628));
  DFFHQX1 \mem_wstrb_reg[3] (.CK (clk), .D (n_9081), .Q (n_5629));
  DFFHQX1 \pcpi_insn_reg[0] (.CK (clk), .D (n_1022), .Q (n_5585));
  DFFHQX1 \pcpi_insn_reg[1] (.CK (clk), .D (n_1021), .Q (n_5586));
  DFFHQX1 \pcpi_insn_reg[2] (.CK (clk), .D (n_998), .Q (n_5587));
  DFFHQX1 \pcpi_insn_reg[3] (.CK (clk), .D (n_1020), .Q (n_5588));
  DFFHQX1 \pcpi_insn_reg[4] (.CK (clk), .D (n_999), .Q (n_5589));
  DFFHQX1 \pcpi_insn_reg[5] (.CK (clk), .D (n_1019), .Q (n_5590));
  DFFHQX1 \pcpi_insn_reg[6] (.CK (clk), .D (n_1018), .Q (n_5591));
  DFFHQX1 \pcpi_insn_reg[7] (.CK (clk), .D (n_1017), .Q (n_5592));
  DFFHQX1 \pcpi_insn_reg[8] (.CK (clk), .D (n_1023), .Q (n_5593));
  DFFHQX1 \pcpi_insn_reg[9] (.CK (clk), .D (n_1016), .Q (n_5594));
  DFFHQX1 \pcpi_insn_reg[10] (.CK (clk), .D (n_1024), .Q (n_5595));
  DFFHQX1 \pcpi_insn_reg[11] (.CK (clk), .D (n_1015), .Q (n_5596));
  DFFHQX1 \pcpi_insn_reg[12] (.CK (clk), .D (n_1025), .Q (n_5597));
  DFFHQX1 \pcpi_insn_reg[13] (.CK (clk), .D (n_1014), .Q (n_5598));
  DFFHQX1 \pcpi_insn_reg[14] (.CK (clk), .D (n_1013), .Q (n_5599));
  DFFHQX1 \pcpi_insn_reg[15] (.CK (clk), .D (n_1012), .Q (n_5600));
  DFFHQX1 \pcpi_insn_reg[16] (.CK (clk), .D (n_995), .Q (n_5601));
  DFFHQX1 \pcpi_insn_reg[17] (.CK (clk), .D (n_1011), .Q (n_5602));
  DFFHQX1 \pcpi_insn_reg[18] (.CK (clk), .D (n_1010), .Q (n_5603));
  DFFHQX1 \pcpi_insn_reg[19] (.CK (clk), .D (n_1009), .Q (n_5604));
  DFFHQX1 \pcpi_insn_reg[20] (.CK (clk), .D (n_1000), .Q (n_5605));
  DFFHQX1 \pcpi_insn_reg[21] (.CK (clk), .D (n_1008), .Q (n_5606));
  DFFHQX1 \pcpi_insn_reg[22] (.CK (clk), .D (n_1007), .Q (n_5607));
  DFFHQX1 \pcpi_insn_reg[23] (.CK (clk), .D (n_1006), .Q (n_5608));
  DFFHQX1 \pcpi_insn_reg[24] (.CK (clk), .D (n_996), .Q (n_5609));
  DFFHQX1 \pcpi_insn_reg[25] (.CK (clk), .D (n_1005), .Q (n_5610));
  DFFHQX1 \pcpi_insn_reg[26] (.CK (clk), .D (n_997), .Q (n_5611));
  DFFHQX1 \pcpi_insn_reg[27] (.CK (clk), .D (n_1004), .Q (n_5612));
  DFFHQX1 \pcpi_insn_reg[28] (.CK (clk), .D (n_1026), .Q (n_5613));
  DFFHQX1 \pcpi_insn_reg[29] (.CK (clk), .D (n_1003), .Q (n_5614));
  DFFHQX1 \pcpi_insn_reg[30] (.CK (clk), .D (n_1002), .Q (n_5615));
  DFFHQX1 \pcpi_insn_reg[31] (.CK (clk), .D (n_1001), .Q (n_5616));
  DFFHQX1 \pcpi_timeout_counter_reg[0] (.CK (clk), .D (n_1540), .Q
       (pcpi_timeout_counter[0]));
  DFFHQX1 \pcpi_timeout_counter_reg[1] (.CK (clk), .D (n_1919), .Q
       (pcpi_timeout_counter[1]));
  DFFHQX1 \pcpi_timeout_counter_reg[2] (.CK (clk), .D (n_1920), .Q
       (pcpi_timeout_counter[2]));
  DFFHQX1 \pcpi_timeout_counter_reg[3] (.CK (clk), .D (n_1553), .Q
       (pcpi_timeout_counter[3]));
  DFFHQX1 pcpi_valid_reg(.CK (clk), .D (n_2295), .Q (n_5617));
  DFFHQX1 prefetched_high_word_reg(.CK (clk), .D (n_2589), .Q
       (prefetched_high_word));
  DFFHQX1 \reg_next_pc_reg[1] (.CK (clk), .D (n_2257), .Q
       (reg_next_pc[1]));
  DFFHQX1 \reg_next_pc_reg[2] (.CK (clk), .D (n_2256), .Q
       (reg_next_pc[2]));
  DFFHQX1 \reg_next_pc_reg[3] (.CK (clk), .D (n_2255), .Q
       (reg_next_pc[3]));
  DFFHQX1 \reg_next_pc_reg[4] (.CK (clk), .D (n_2254), .Q
       (reg_next_pc[4]));
  DFFHQX1 \reg_next_pc_reg[5] (.CK (clk), .D (n_2253), .Q
       (reg_next_pc[5]));
  DFFHQX1 \reg_next_pc_reg[6] (.CK (clk), .D (n_2252), .Q
       (reg_next_pc[6]));
  DFFHQX1 \reg_next_pc_reg[7] (.CK (clk), .D (n_2251), .Q
       (reg_next_pc[7]));
  DFFHQX1 \reg_next_pc_reg[8] (.CK (clk), .D (n_2250), .Q
       (reg_next_pc[8]));
  DFFHQX1 \reg_next_pc_reg[9] (.CK (clk), .D (n_2249), .Q
       (reg_next_pc[9]));
  DFFHQX1 \reg_next_pc_reg[10] (.CK (clk), .D (n_2248), .Q
       (reg_next_pc[10]));
  DFFHQX1 \reg_next_pc_reg[11] (.CK (clk), .D (n_2247), .Q
       (reg_next_pc[11]));
  DFFHQX1 \reg_next_pc_reg[12] (.CK (clk), .D (n_2246), .Q
       (reg_next_pc[12]));
  DFFHQX1 \reg_next_pc_reg[13] (.CK (clk), .D (n_2245), .Q
       (reg_next_pc[13]));
  DFFHQX1 \reg_next_pc_reg[14] (.CK (clk), .D (n_2244), .Q
       (reg_next_pc[14]));
  DFFHQX1 \reg_next_pc_reg[15] (.CK (clk), .D (n_2243), .Q
       (reg_next_pc[15]));
  DFFHQX1 \reg_next_pc_reg[16] (.CK (clk), .D (n_2242), .Q
       (reg_next_pc[16]));
  DFFHQX1 \reg_next_pc_reg[17] (.CK (clk), .D (n_2241), .Q
       (reg_next_pc[17]));
  DFFHQX1 \reg_next_pc_reg[18] (.CK (clk), .D (n_2240), .Q
       (reg_next_pc[18]));
  DFFHQX1 \reg_next_pc_reg[19] (.CK (clk), .D (n_2225), .Q
       (reg_next_pc[19]));
  DFFHQX1 \reg_next_pc_reg[20] (.CK (clk), .D (n_2239), .Q
       (reg_next_pc[20]));
  DFFHQX1 \reg_next_pc_reg[21] (.CK (clk), .D (n_2238), .Q
       (reg_next_pc[21]));
  DFFHQX1 \reg_next_pc_reg[22] (.CK (clk), .D (n_2237), .Q
       (reg_next_pc[22]));
  DFFHQX1 \reg_next_pc_reg[23] (.CK (clk), .D (n_2236), .Q
       (reg_next_pc[23]));
  DFFHQX1 \reg_next_pc_reg[24] (.CK (clk), .D (n_2235), .Q
       (reg_next_pc[24]));
  DFFHQX1 \reg_next_pc_reg[25] (.CK (clk), .D (n_2234), .Q
       (reg_next_pc[25]));
  DFFHQX1 \reg_next_pc_reg[26] (.CK (clk), .D (n_2226), .Q
       (reg_next_pc[26]));
  DFFHQX1 \reg_next_pc_reg[27] (.CK (clk), .D (n_2233), .Q
       (reg_next_pc[27]));
  DFFHQX1 \reg_next_pc_reg[28] (.CK (clk), .D (n_2232), .Q
       (reg_next_pc[28]));
  DFFHQX1 \reg_next_pc_reg[29] (.CK (clk), .D (n_2231), .Q
       (reg_next_pc[29]));
  DFFHQX1 \reg_next_pc_reg[30] (.CK (clk), .D (n_2230), .Q
       (reg_next_pc[30]));
  DFFHQX1 \reg_next_pc_reg[31] (.CK (clk), .D (n_2227), .Q
       (reg_next_pc[31]));
  DFFHQX1 \reg_op1_reg[0] (.CK (clk), .D (n_5234), .Q (reg_op1[0]));
  DFFHQX1 \reg_op1_reg[1] (.CK (clk), .D (n_5231), .Q (\reg_op1[1]_9638
       ));
  DFFHQX1 \reg_op1_reg[2] (.CK (clk), .D (n_5160), .Q (\reg_op1[2]_9639
       ));
  DFFHQX1 \reg_op1_reg[3] (.CK (clk), .D (n_5161), .Q (\reg_op1[3]_9640
       ));
  DFFHQX1 \reg_op1_reg[4] (.CK (clk), .D (n_5255), .Q (\reg_op1[4]_9641
       ));
  DFFHQX1 \reg_op1_reg[5] (.CK (clk), .D (n_5252), .Q (\reg_op1[5]_9642
       ));
  DFFHQX1 \reg_op1_reg[6] (.CK (clk), .D (n_5237), .Q (\reg_op1[6]_9643
       ));
  DFFHQX1 \reg_op1_reg[7] (.CK (clk), .D (n_5243), .Q (\reg_op1[7]_9644
       ));
  DFFHQX1 \reg_op1_reg[8] (.CK (clk), .D (n_5253), .Q (\reg_op1[8]_9645
       ));
  DFFHQX1 \reg_op1_reg[9] (.CK (clk), .D (n_5254), .Q (\reg_op1[9]_9646
       ));
  DFFHQX1 \reg_op1_reg[10] (.CK (clk), .D (n_5246), .Q
       (\reg_op1[10]_9647 ));
  DFFHQX1 \reg_op1_reg[11] (.CK (clk), .D (n_5250), .Q
       (\reg_op1[11]_9648 ));
  DFFHQX1 \reg_op1_reg[12] (.CK (clk), .D (n_5249), .Q
       (\reg_op1[12]_9649 ));
  DFFHQX1 \reg_op1_reg[13] (.CK (clk), .D (n_5248), .Q
       (\reg_op1[13]_9650 ));
  DFFHQX1 \reg_op1_reg[14] (.CK (clk), .D (n_5176), .Q
       (\reg_op1[14]_9651 ));
  DFFHQX1 \reg_op1_reg[15] (.CK (clk), .D (n_5238), .Q
       (\reg_op1[15]_9652 ));
  DFFHQX1 \reg_op1_reg[16] (.CK (clk), .D (n_5175), .Q
       (\reg_op1[16]_9653 ));
  DFFHQX1 \reg_op1_reg[17] (.CK (clk), .D (n_5247), .Q
       (\reg_op1[17]_9654 ));
  DFFHQX1 \reg_op1_reg[18] (.CK (clk), .D (n_5214), .Q
       (\reg_op1[18]_9655 ));
  DFFHQX1 \reg_op1_reg[19] (.CK (clk), .D (n_5233), .Q
       (\reg_op1[19]_9656 ));
  DFFHQX1 \reg_op1_reg[20] (.CK (clk), .D (n_5206), .Q
       (\reg_op1[20]_9657 ));
  DFFHQX1 \reg_op1_reg[21] (.CK (clk), .D (n_5204), .Q
       (\reg_op1[21]_9658 ));
  DFFHQX1 \reg_op1_reg[22] (.CK (clk), .D (n_5232), .Q
       (\reg_op1[22]_9659 ));
  DFFHQX1 \reg_op1_reg[23] (.CK (clk), .D (n_5241), .Q
       (\reg_op1[23]_9660 ));
  DFFHQX1 \reg_op1_reg[24] (.CK (clk), .D (n_5251), .Q
       (\reg_op1[24]_9661 ));
  DFFHQX1 \reg_op1_reg[25] (.CK (clk), .D (n_5174), .Q
       (\reg_op1[25]_9662 ));
  DFFHQX1 \reg_op1_reg[26] (.CK (clk), .D (n_5245), .Q
       (\reg_op1[26]_9663 ));
  DFFHQX1 \reg_op1_reg[27] (.CK (clk), .D (n_5244), .Q
       (\reg_op1[27]_9664 ));
  DFFHQX1 \reg_op1_reg[28] (.CK (clk), .D (n_5242), .Q
       (\reg_op1[28]_9665 ));
  DFFHQX1 \reg_op1_reg[29] (.CK (clk), .D (n_5256), .Q
       (\reg_op1[29]_9666 ));
  DFFHQX1 \reg_op1_reg[30] (.CK (clk), .D (n_5179), .Q
       (\reg_op1[30]_9667 ));
  DFFHQX1 \reg_op1_reg[31] (.CK (clk), .D (n_5180), .Q
       (\reg_op1[31]_9668 ));
  DFFHQX1 \reg_op2_reg[0] (.CK (clk), .D (n_4852), .Q (\reg_op2[0]_9669
       ));
  DFFHQX1 \reg_op2_reg[1] (.CK (clk), .D (n_4851), .Q (\reg_op2[1]_9670
       ));
  DFFHQX1 \reg_op2_reg[2] (.CK (clk), .D (n_4528), .Q (\reg_op2[2]_9671
       ));
  DFFHQX1 \reg_op2_reg[3] (.CK (clk), .D (n_4527), .Q (\reg_op2[3]_9672
       ));
  DFFHQX1 \reg_op2_reg[4] (.CK (clk), .D (n_4850), .Q (\reg_op2[4]_9673
       ));
  DFFHQX1 \reg_op2_reg[5] (.CK (clk), .D (n_4765), .Q (\reg_op2[5]_9674
       ));
  DFFHQX1 \reg_op2_reg[6] (.CK (clk), .D (n_4764), .Q (\reg_op2[6]_9675
       ));
  DFFHQX1 \reg_op2_reg[7] (.CK (clk), .D (n_4973), .Q (\reg_op2[7]_9676
       ));
  DFFHQX1 \reg_op2_reg[8] (.CK (clk), .D (n_4970), .Q (\reg_op2[8]_9677
       ));
  DFFHQX1 \reg_op2_reg[9] (.CK (clk), .D (n_4969), .Q (\reg_op2[9]_9678
       ));
  DFFHQX1 \reg_op2_reg[10] (.CK (clk), .D (n_4763), .Q
       (\reg_op2[10]_9679 ));
  DFFHQX1 \reg_op2_reg[11] (.CK (clk), .D (n_4968), .Q
       (\reg_op2[11]_9680 ));
  DFFHQX1 \reg_op2_reg[12] (.CK (clk), .D (n_4967), .Q
       (\reg_op2[12]_9681 ));
  DFFHQX1 \reg_op2_reg[13] (.CK (clk), .D (n_4966), .Q
       (\reg_op2[13]_9682 ));
  DFFHQX1 \reg_op2_reg[14] (.CK (clk), .D (n_4965), .Q
       (\reg_op2[14]_9683 ));
  DFFHQX1 \reg_op2_reg[15] (.CK (clk), .D (n_4964), .Q
       (\reg_op2[15]_9684 ));
  DFFHQX1 \reg_op2_reg[16] (.CK (clk), .D (n_4963), .Q
       (\reg_op2[16]_9685 ));
  DFFHQX1 \reg_op2_reg[17] (.CK (clk), .D (n_4762), .Q
       (\reg_op2[17]_9686 ));
  DFFHQX1 \reg_op2_reg[18] (.CK (clk), .D (n_4960), .Q
       (\reg_op2[18]_9687 ));
  DFFHQX1 \reg_op2_reg[19] (.CK (clk), .D (n_4971), .Q
       (\reg_op2[19]_9688 ));
  DFFHQX1 \reg_op2_reg[20] (.CK (clk), .D (n_4961), .Q
       (\reg_op2[20]_9689 ));
  DFFHQX1 \reg_op2_reg[21] (.CK (clk), .D (n_4959), .Q
       (\reg_op2[21]_9690 ));
  DFFHQX1 \reg_op2_reg[22] (.CK (clk), .D (n_4958), .Q
       (\reg_op2[22]_9691 ));
  DFFHQX1 \reg_op2_reg[23] (.CK (clk), .D (n_4761), .Q
       (\reg_op2[23]_9692 ));
  DFFHQX1 \reg_op2_reg[24] (.CK (clk), .D (n_4972), .Q
       (\reg_op2[24]_9693 ));
  DFFHQX1 \reg_op2_reg[25] (.CK (clk), .D (n_4957), .Q
       (\reg_op2[25]_9694 ));
  DFFHQX1 \reg_op2_reg[26] (.CK (clk), .D (n_4760), .Q
       (\reg_op2[26]_9695 ));
  DFFHQX1 \reg_op2_reg[27] (.CK (clk), .D (n_4956), .Q
       (\reg_op2[27]_9696 ));
  DFFHQX1 \reg_op2_reg[28] (.CK (clk), .D (n_4759), .Q
       (\reg_op2[28]_9697 ));
  DFFHQX1 \reg_op2_reg[29] (.CK (clk), .D (n_4978), .Q
       (\reg_op2[29]_9698 ));
  DFFHQX1 \reg_op2_reg[30] (.CK (clk), .D (n_4955), .Q
       (\reg_op2[30]_9699 ));
  DFFHQX1 \reg_op2_reg[31] (.CK (clk), .D (n_4954), .Q
       (\reg_op2[31]_9700 ));
  DFFHQX1 \reg_out_reg[1] (.CK (clk), .D (n_2474), .Q (reg_out[1]));
  DFFHQX1 \reg_out_reg[2] (.CK (clk), .D (n_2450), .Q (reg_out[2]));
  DFFHQX1 \reg_out_reg[3] (.CK (clk), .D (n_2454), .Q (reg_out[3]));
  DFFHQX1 \reg_out_reg[4] (.CK (clk), .D (n_2466), .Q (reg_out[4]));
  DFFHQX1 \reg_out_reg[5] (.CK (clk), .D (n_2467), .Q (reg_out[5]));
  DFFHQX1 \reg_out_reg[6] (.CK (clk), .D (n_2468), .Q (reg_out[6]));
  DFFHQX1 \reg_out_reg[7] (.CK (clk), .D (n_2371), .Q (reg_out[7]));
  DFFHQX1 \reg_out_reg[8] (.CK (clk), .D (n_2582), .Q (reg_out[8]));
  DFFHQX1 \reg_out_reg[9] (.CK (clk), .D (n_2559), .Q (reg_out[9]));
  DFFHQX1 \reg_out_reg[10] (.CK (clk), .D (n_2581), .Q (reg_out[10]));
  DFFHQX1 \reg_out_reg[11] (.CK (clk), .D (n_2580), .Q (reg_out[11]));
  DFFHQX1 \reg_out_reg[12] (.CK (clk), .D (n_2579), .Q (reg_out[12]));
  DFFHQX1 \reg_out_reg[13] (.CK (clk), .D (n_2578), .Q (reg_out[13]));
  DFFHQX1 \reg_out_reg[14] (.CK (clk), .D (n_2577), .Q (reg_out[14]));
  DFFHQX1 \reg_out_reg[15] (.CK (clk), .D (n_2469), .Q (reg_out[15]));
  DFFHQX1 \reg_out_reg[16] (.CK (clk), .D (n_2488), .Q (reg_out[16]));
  DFFHQX1 \reg_out_reg[17] (.CK (clk), .D (n_2455), .Q (reg_out[17]));
  DFFHQX1 \reg_out_reg[18] (.CK (clk), .D (n_2453), .Q (reg_out[18]));
  DFFHQX1 \reg_out_reg[19] (.CK (clk), .D (n_2452), .Q (reg_out[19]));
  DFFHQX1 \reg_out_reg[20] (.CK (clk), .D (n_2451), .Q (reg_out[20]));
  DFFHQX1 \reg_out_reg[21] (.CK (clk), .D (n_2465), .Q (reg_out[21]));
  DFFHQX1 \reg_out_reg[22] (.CK (clk), .D (n_2464), .Q (reg_out[22]));
  DFFHQX1 \reg_out_reg[23] (.CK (clk), .D (n_2463), .Q (reg_out[23]));
  DFFHQX1 \reg_out_reg[24] (.CK (clk), .D (n_2462), .Q (reg_out[24]));
  DFFHQX1 \reg_out_reg[25] (.CK (clk), .D (n_2461), .Q (reg_out[25]));
  DFFHQX1 \reg_out_reg[26] (.CK (clk), .D (n_2460), .Q (reg_out[26]));
  DFFHQX1 \reg_out_reg[27] (.CK (clk), .D (n_2459), .Q (reg_out[27]));
  DFFHQX1 \reg_out_reg[28] (.CK (clk), .D (n_2458), .Q (reg_out[28]));
  DFFHQX1 \reg_out_reg[29] (.CK (clk), .D (n_2457), .Q (reg_out[29]));
  DFFHQX1 \reg_out_reg[30] (.CK (clk), .D (n_2456), .Q (reg_out[30]));
  DFFHQX1 \reg_out_reg[31] (.CK (clk), .D (n_3411), .Q (reg_out[31]));
  DFFHQX1 \reg_pc_reg[1] (.CK (clk), .D (n_11826), .Q (reg_pc[1]));
  DFFHQX1 \reg_pc_reg[2] (.CK (clk), .D (n_11821), .Q (reg_pc[2]));
  DFFHQX1 \reg_pc_reg[3] (.CK (clk), .D (n_11825), .Q (reg_pc[3]));
  DFFHQX1 \reg_pc_reg[4] (.CK (clk), .D (n_11823), .Q (reg_pc[4]));
  DFFHQX1 \reg_pc_reg[5] (.CK (clk), .D (n_11822), .Q (reg_pc[5]));
  DFFHQX1 \reg_pc_reg[6] (.CK (clk), .D (n_11824), .Q (reg_pc[6]));
  DFFHQX1 \reg_pc_reg[7] (.CK (clk), .D (n_11831), .Q (reg_pc[7]));
  DFFHQX1 \reg_pc_reg[8] (.CK (clk), .D (n_11803), .Q (reg_pc[8]));
  DFFHQX1 \reg_pc_reg[9] (.CK (clk), .D (n_11802), .Q (reg_pc[9]));
  DFFHQX1 \reg_pc_reg[10] (.CK (clk), .D (n_11820), .Q (reg_pc[10]));
  DFFHQX1 \reg_pc_reg[11] (.CK (clk), .D (n_11827), .Q (reg_pc[11]));
  DFFHQX1 \reg_pc_reg[12] (.CK (clk), .D (n_11812), .Q (reg_pc[12]));
  DFFHQX1 \reg_pc_reg[13] (.CK (clk), .D (n_11817), .Q (reg_pc[13]));
  DFFHQX1 \reg_pc_reg[14] (.CK (clk), .D (n_11814), .Q (reg_pc[14]));
  DFFHQX1 \reg_pc_reg[15] (.CK (clk), .D (n_11807), .Q (reg_pc[15]));
  DFFHQX1 \reg_pc_reg[16] (.CK (clk), .D (n_11801), .Q (reg_pc[16]));
  DFFHQX1 \reg_pc_reg[17] (.CK (clk), .D (n_11805), .Q (reg_pc[17]));
  DFFHQX1 \reg_pc_reg[18] (.CK (clk), .D (n_11819), .Q (reg_pc[18]));
  DFFHQX1 \reg_pc_reg[19] (.CK (clk), .D (n_11809), .Q (reg_pc[19]));
  DFFHQX1 \reg_pc_reg[20] (.CK (clk), .D (n_11810), .Q (reg_pc[20]));
  DFFHQX1 \reg_pc_reg[21] (.CK (clk), .D (n_11813), .Q (reg_pc[21]));
  DFFHQX1 \reg_pc_reg[22] (.CK (clk), .D (n_11830), .Q (reg_pc[22]));
  DFFHQX1 \reg_pc_reg[23] (.CK (clk), .D (n_11816), .Q (reg_pc[23]));
  DFFHQX1 \reg_pc_reg[24] (.CK (clk), .D (n_11806), .Q (reg_pc[24]));
  DFFHQX1 \reg_pc_reg[25] (.CK (clk), .D (n_11804), .Q (reg_pc[25]));
  DFFHQX1 \reg_pc_reg[26] (.CK (clk), .D (n_11828), .Q (reg_pc[26]));
  DFFHQX1 \reg_pc_reg[27] (.CK (clk), .D (n_11818), .Q (reg_pc[27]));
  DFFHQX1 \reg_pc_reg[28] (.CK (clk), .D (n_11808), .Q (reg_pc[28]));
  DFFHQX1 \reg_pc_reg[29] (.CK (clk), .D (n_11811), .Q (reg_pc[29]));
  DFFHQX1 \reg_pc_reg[30] (.CK (clk), .D (n_11829), .Q (reg_pc[30]));
  DFFHQX1 \reg_pc_reg[31] (.CK (clk), .D (n_11815), .Q (reg_pc[31]));
  DFFHQX1 \reg_sh_reg[0] (.CK (clk), .D (n_4854), .Q (reg_sh[0]));
  DFFHQX1 \reg_sh_reg[1] (.CK (clk), .D (n_4919), .Q (reg_sh[1]));
  DFFHQX1 \reg_sh_reg[2] (.CK (clk), .D (n_4708), .Q (reg_sh[2]));
  DFFHQX1 \reg_sh_reg[3] (.CK (clk), .D (n_3470), .Q (reg_sh[3]));
  DFFHQX1 \reg_sh_reg[4] (.CK (clk), .D (n_4906), .Q (reg_sh[4]));
  DFFHQX1 trap_reg(.CK (clk), .D (n_890), .Q (n_5693));
  OAI21X1 g174701__7098(.A0 (n_953), .A1 (n_5521), .B0 (n_1361), .Y
       (n_5528));
  NOR2X1 g174703__6131(.A (n_544), .B (n_5525), .Y (n_5527));
  NOR2X1 g174704__1881(.A (n_544), .B (n_5524), .Y (n_5526));
  AOI21X1 g174705__5115(.A0 (latched_store), .A1 (n_2512), .B0
       (n_5522), .Y (n_5525));
  MX2X1 g174706__7482(.A (n_5517), .B (n_555), .S0 (n_779), .Y
       (n_5524));
  MX2X1 g174707__4733(.A (n_5516), .B (n_4710), .S0 (n_5520), .Y
       (n_5523));
  NOR2X1 g174708__6161(.A (n_2512), .B (n_5519), .Y (n_5522));
  NOR2X1 g174709__9315(.A (cpu_state[5]), .B (n_5518), .Y (n_5521));
  NOR2X1 g174711__9945(.A (n_850), .B (n_5516), .Y (n_5520));
  AOI221X1 g174712__2883(.A0 (n_2388), .A1 (n_5511), .B0
       (cpu_state[5]), .B1 (n_297), .C0 (n_852), .Y (n_5519));
  OAI211X1 g174713__2346(.A0 (n_613), .A1 (n_5512), .B0 (n_615), .C0
       (n_11), .Y (n_5518));
  AOI221X1 g174714__1666(.A0 (instr_jalr), .A1 (n_849), .B0
       (instr_jal), .B1 (n_666), .C0 (n_5514), .Y (n_5517));
  AND2X1 g174715__7410(.A (n_5514), .B (n_543), .Y (n_5516));
  NAND4XL g174716__6417(.A (n_1263), .B (n_1916), .C (n_1267), .D
       (n_5513), .Y (n_5515));
  AND2X1 g174717__5477(.A (n_5512), .B (cpu_state[3]), .Y (n_5514));
  AOI22XL g174718__2398(.A0 (is_compare), .A1 (n_5510), .B0
       (is_lui_auipc_jal_jalr_addi_add_sub), .B1 (n_6625), .Y (n_5513));
  AND2X1 g174719__5107(.A (n_5510), .B (is_beq_bne_blt_bge_bltu_bgeu),
       .Y (n_5512));
  NAND2BX1 g174720__6260(.AN (n_5510), .B
       (is_beq_bne_blt_bge_bltu_bgeu), .Y (n_5511));
  NAND3X1 g174721__4319(.A (n_5508), .B (n_5509), .C (n_5507), .Y
       (n_5510));
  AOI22X1 g174722__8428(.A0 (instr_bgeu), .A1 (n_5506), .B0
       (instr_bne), .B1 (n_5030), .Y (n_5509));
  AOI22XL g174723__5526(.A0 (is_slti_blt_slt), .A1 (n_5504), .B0
       (instr_beq), .B1 (n_5029), .Y (n_5508));
  AOI22XL g174724__6783(.A0 (is_sltiu_bltu_sltu), .A1 (n_5505), .B0
       (instr_bge), .B1 (n_5503), .Y (n_5507));
  INVX1 g174725(.A (n_5505), .Y (n_5506));
  AOI21X1 g174726__3680(.A0 (n_868), .A1 (n_5501), .B0 (n_866), .Y
       (n_5505));
  INVX1 g174727(.A (n_5503), .Y (n_5504));
  NAND2X1 g174728__1617(.A (n_868), .B (n_5502), .Y (n_5503));
  NAND2BX1 g174729__2802(.AN (n_866), .B (n_5501), .Y (n_5502));
  OAI2BB1X1 g174730__1705(.A0N (n_6552), .A1N (n_5500), .B0 (n_6553),
       .Y (n_5501));
  OAI22X1 g174731__5122(.A0 (n_816), .A1 (n_5499), .B0
       (\reg_op2[29]_9698 ), .B1 (n_716), .Y (n_5500));
  AOI22X1 g174732__8246(.A0 (\genblk2.pcpi_div_minus_2470_59_n_479 ),
       .A1 (n_5483), .B0 (\reg_op1[28]_9665 ), .B1 (n_5465), .Y
       (n_5499));
  OAI2BB1X1 g174765__7098(.A0N (\genblk2.pcpi_div_dividend [14]), .A1N
       (n_5270), .B0 (n_5464), .Y (n_5498));
  OAI2BB1X1 g174766__6131(.A0N (\genblk2.pcpi_div_dividend [0]), .A1N
       (n_5270), .B0 (n_5463), .Y (n_5497));
  OAI2BB1X1 g174767__1881(.A0N (\genblk2.pcpi_div_dividend [1]), .A1N
       (n_5270), .B0 (n_5462), .Y (n_5496));
  OAI2BB1X1 g174768__5115(.A0N (\genblk2.pcpi_div_dividend [2]), .A1N
       (n_5270), .B0 (n_5461), .Y (n_5495));
  OAI2BB1X1 g174769__7482(.A0N (\genblk2.pcpi_div_dividend [3]), .A1N
       (n_5270), .B0 (n_5460), .Y (n_5494));
  OAI2BB1X1 g174770__4733(.A0N (\genblk2.pcpi_div_dividend [5]), .A1N
       (n_5270), .B0 (n_5458), .Y (n_5493));
  OAI2BB1X1 g174771__6161(.A0N (\genblk2.pcpi_div_dividend [4]), .A1N
       (n_5270), .B0 (n_5459), .Y (n_5492));
  OAI2BB1X1 g174772__9315(.A0N (\genblk2.pcpi_div_dividend [6]), .A1N
       (n_5270), .B0 (n_5457), .Y (n_5491));
  OAI2BB1X1 g174773__9945(.A0N (\genblk2.pcpi_div_dividend [7]), .A1N
       (n_5270), .B0 (n_5456), .Y (n_5490));
  OAI2BB1X1 g174774__2883(.A0N (\genblk2.pcpi_div_dividend [8]), .A1N
       (n_5270), .B0 (n_5455), .Y (n_5489));
  OAI2BB1X1 g174775__2346(.A0N (\genblk2.pcpi_div_dividend [10]), .A1N
       (n_5270), .B0 (n_5453), .Y (n_5488));
  OAI2BB1X1 g174776__1666(.A0N (\genblk2.pcpi_div_dividend [9]), .A1N
       (n_5270), .B0 (n_5454), .Y (n_5487));
  OAI2BB1X1 g174777__7410(.A0N (\genblk2.pcpi_div_dividend [11]), .A1N
       (n_5270), .B0 (n_5452), .Y (n_5486));
  OAI2BB1X1 g174778__6417(.A0N (\genblk2.pcpi_div_dividend [12]), .A1N
       (n_5270), .B0 (n_5451), .Y (n_5485));
  OAI2BB1X1 g174779__5477(.A0N (\genblk2.pcpi_div_dividend [13]), .A1N
       (n_5270), .B0 (n_5450), .Y (n_5484));
  OR2X1 g174780__2398(.A (\reg_op1[28]_9665 ), .B (n_5465), .Y
       (n_5483));
  OAI2BB1X1 g174781__5107(.A0N (\genblk2.pcpi_div_dividend [15]), .A1N
       (n_5270), .B0 (n_5449), .Y (n_5482));
  OAI2BB1X1 g174782__6260(.A0N (\genblk2.pcpi_div_dividend [16]), .A1N
       (n_5270), .B0 (n_5448), .Y (n_5481));
  OAI2BB1X1 g174783__4319(.A0N (\genblk2.pcpi_div_dividend [17]), .A1N
       (n_5270), .B0 (n_5447), .Y (n_5480));
  OAI2BB1X1 g174784__8428(.A0N (\genblk2.pcpi_div_dividend [18]), .A1N
       (n_5270), .B0 (n_5446), .Y (n_5479));
  OAI2BB1X1 g174785__5526(.A0N (\genblk2.pcpi_div_dividend [19]), .A1N
       (n_5270), .B0 (n_5445), .Y (n_5478));
  OAI2BB1X1 g174786__6783(.A0N (\genblk2.pcpi_div_dividend [22]), .A1N
       (n_5270), .B0 (n_5442), .Y (n_5477));
  OAI2BB1X1 g174787__3680(.A0N (\genblk2.pcpi_div_dividend [20]), .A1N
       (n_5270), .B0 (n_5444), .Y (n_5476));
  OAI2BB1X1 g174788__1617(.A0N (\genblk2.pcpi_div_dividend [23]), .A1N
       (n_5270), .B0 (n_5441), .Y (n_5475));
  OAI2BB1X1 g174789__2802(.A0N (\genblk2.pcpi_div_dividend [21]), .A1N
       (n_5270), .B0 (n_5443), .Y (n_5474));
  OAI2BB1X1 g174790__1705(.A0N (\genblk2.pcpi_div_dividend [24]), .A1N
       (n_5270), .B0 (n_5440), .Y (n_5473));
  OAI2BB1X1 g174791__5122(.A0N (\genblk2.pcpi_div_dividend [25]), .A1N
       (n_5270), .B0 (n_5439), .Y (n_5472));
  OAI2BB1X1 g174792__8246(.A0N (\genblk2.pcpi_div_dividend [26]), .A1N
       (n_5270), .B0 (n_5438), .Y (n_5471));
  OAI2BB1X1 g174793__7098(.A0N (\genblk2.pcpi_div_dividend [27]), .A1N
       (n_5270), .B0 (n_5437), .Y (n_5470));
  OAI2BB1X1 g174794__6131(.A0N (\genblk2.pcpi_div_dividend [28]), .A1N
       (n_5270), .B0 (n_5436), .Y (n_5469));
  OAI2BB1X1 g174795__1881(.A0N (\genblk2.pcpi_div_dividend [29]), .A1N
       (n_5270), .B0 (n_5435), .Y (n_5468));
  OAI2BB1X1 g174796__5115(.A0N (\genblk2.pcpi_div_dividend [30]), .A1N
       (n_5270), .B0 (n_5433), .Y (n_5467));
  OAI2BB1X1 g174797__7482(.A0N (\genblk2.pcpi_div_dividend [31]), .A1N
       (n_5270), .B0 (n_5434), .Y (n_5466));
  AOI22XL g174798__4733(.A0 (\genblk2.pcpi_div_n_1947 ), .A1 (n_5431),
       .B0 (\reg_op1[14]_9651 ), .B1 (n_460), .Y (n_5464));
  AOI22XL g174799__6161(.A0 (\genblk2.pcpi_div_n_1961 ), .A1 (n_5431),
       .B0 (reg_op1[0]), .B1 (n_460), .Y (n_5463));
  AOI22XL g174800__9315(.A0 (\genblk2.pcpi_div_n_1960 ), .A1 (n_5431),
       .B0 (\reg_op1[1]_9638 ), .B1 (n_460), .Y (n_5462));
  AOI22XL g174801__9945(.A0 (\genblk2.pcpi_div_n_1959 ), .A1 (n_5431),
       .B0 (\reg_op1[2]_9639 ), .B1 (n_460), .Y (n_5461));
  AOI22XL g174802__2883(.A0 (\genblk2.pcpi_div_n_1958 ), .A1 (n_5431),
       .B0 (\reg_op1[3]_9640 ), .B1 (n_460), .Y (n_5460));
  AOI22XL g174803__2346(.A0 (\genblk2.pcpi_div_n_1957 ), .A1 (n_5431),
       .B0 (\reg_op1[4]_9641 ), .B1 (n_460), .Y (n_5459));
  AOI22XL g174804__1666(.A0 (\genblk2.pcpi_div_n_1956 ), .A1 (n_5431),
       .B0 (\reg_op1[5]_9642 ), .B1 (n_460), .Y (n_5458));
  AOI22XL g174805__7410(.A0 (\genblk2.pcpi_div_n_1955 ), .A1 (n_5431),
       .B0 (\reg_op1[6]_9643 ), .B1 (n_460), .Y (n_5457));
  AOI22XL g174806__6417(.A0 (\genblk2.pcpi_div_n_1954 ), .A1 (n_5431),
       .B0 (\reg_op1[7]_9644 ), .B1 (n_460), .Y (n_5456));
  AOI22XL g174807__5477(.A0 (\genblk2.pcpi_div_n_1953 ), .A1 (n_5431),
       .B0 (\reg_op1[8]_9645 ), .B1 (n_460), .Y (n_5455));
  AOI22XL g174808__2398(.A0 (\genblk2.pcpi_div_n_1952 ), .A1 (n_5431),
       .B0 (\reg_op1[9]_9646 ), .B1 (n_460), .Y (n_5454));
  AOI22XL g174809__5107(.A0 (\genblk2.pcpi_div_n_1951 ), .A1 (n_5431),
       .B0 (\reg_op1[10]_9647 ), .B1 (n_460), .Y (n_5453));
  AOI22XL g174810__6260(.A0 (\genblk2.pcpi_div_n_1950 ), .A1 (n_5431),
       .B0 (\reg_op1[11]_9648 ), .B1 (n_460), .Y (n_5452));
  AOI22XL g174811__4319(.A0 (\genblk2.pcpi_div_n_1949 ), .A1 (n_5431),
       .B0 (\reg_op1[12]_9649 ), .B1 (n_460), .Y (n_5451));
  AOI22XL g174812__8428(.A0 (\genblk2.pcpi_div_n_1948 ), .A1 (n_5431),
       .B0 (\reg_op1[13]_9650 ), .B1 (n_460), .Y (n_5450));
  OAI211X1 g174813__5526(.A0 (n_876), .A1 (n_1422), .B0 (n_1423), .C0
       (n_5432), .Y (n_5465));
  AOI22XL g174814__6783(.A0 (\genblk2.pcpi_div_n_1946 ), .A1 (n_5431),
       .B0 (\reg_op1[15]_9652 ), .B1 (n_460), .Y (n_5449));
  AOI22XL g174815__3680(.A0 (\genblk2.pcpi_div_n_1945 ), .A1 (n_5431),
       .B0 (\reg_op1[16]_9653 ), .B1 (n_460), .Y (n_5448));
  AOI22XL g174816__1617(.A0 (\genblk2.pcpi_div_n_1944 ), .A1 (n_5431),
       .B0 (\reg_op1[17]_9654 ), .B1 (n_460), .Y (n_5447));
  AOI22XL g174817__2802(.A0 (\genblk2.pcpi_div_n_1943 ), .A1 (n_5431),
       .B0 (\reg_op1[18]_9655 ), .B1 (n_460), .Y (n_5446));
  AOI22XL g174818__1705(.A0 (n_5431), .A1 (\genblk2.pcpi_div_n_1942 ),
       .B0 (\reg_op1[19]_9656 ), .B1 (n_460), .Y (n_5445));
  AOI22XL g174819__5122(.A0 (n_5431), .A1 (\genblk2.pcpi_div_n_1941 ),
       .B0 (\reg_op1[20]_9657 ), .B1 (n_460), .Y (n_5444));
  AOI22XL g174820__8246(.A0 (n_5431), .A1 (\genblk2.pcpi_div_n_1940 ),
       .B0 (\reg_op1[21]_9658 ), .B1 (n_460), .Y (n_5443));
  AOI22XL g174821__7098(.A0 (n_5431), .A1 (\genblk2.pcpi_div_n_1939 ),
       .B0 (\reg_op1[22]_9659 ), .B1 (n_460), .Y (n_5442));
  AOI22XL g174822__6131(.A0 (n_5431), .A1 (\genblk2.pcpi_div_n_1938 ),
       .B0 (\reg_op1[23]_9660 ), .B1 (n_460), .Y (n_5441));
  AOI22XL g174823__1881(.A0 (n_5431), .A1 (\genblk2.pcpi_div_n_1937 ),
       .B0 (\reg_op1[24]_9661 ), .B1 (n_460), .Y (n_5440));
  AOI22XL g174824__5115(.A0 (n_5431), .A1 (\genblk2.pcpi_div_n_1936 ),
       .B0 (\reg_op1[25]_9662 ), .B1 (n_460), .Y (n_5439));
  AOI22XL g174825__7482(.A0 (n_5431), .A1 (\genblk2.pcpi_div_n_1935 ),
       .B0 (\reg_op1[26]_9663 ), .B1 (n_460), .Y (n_5438));
  AOI22XL g174826__4733(.A0 (n_5431), .A1 (\genblk2.pcpi_div_n_1934 ),
       .B0 (\reg_op1[27]_9664 ), .B1 (n_460), .Y (n_5437));
  AOI22XL g174827__6161(.A0 (n_5431), .A1 (\genblk2.pcpi_div_n_1933 ),
       .B0 (\reg_op1[28]_9665 ), .B1 (n_460), .Y (n_5436));
  AOI22XL g174828__9315(.A0 (n_5431), .A1 (\genblk2.pcpi_div_n_1932 ),
       .B0 (\reg_op1[29]_9666 ), .B1 (n_460), .Y (n_5435));
  AOI22XL g174829__9945(.A0 (n_5431), .A1 (\genblk2.pcpi_div_n_1930 ),
       .B0 (\reg_op1[31]_9668 ), .B1 (n_460), .Y (n_5434));
  AOI22XL g174830__2883(.A0 (n_5431), .A1 (\genblk2.pcpi_div_n_1931 ),
       .B0 (\reg_op1[30]_9667 ), .B1 (n_460), .Y (n_5433));
  AOI21X1 g174895__2346(.A0 (n_156), .A1 (n_5267), .B0 (n_778), .Y
       (n_5432));
  NAND2X1 g174961__7410(.A (n_2108), .B (n_5313), .Y (n_5429));
  NAND2X1 g174962__6417(.A (n_2107), .B (n_5312), .Y (n_5428));
  NAND2X1 g174963__5477(.A (n_2106), .B (n_5311), .Y (n_5427));
  NAND2X1 g174964__2398(.A (n_5304), .B (n_2105), .Y (n_5426));
  OAI211X1 g174965__5107(.A0 (n_629), .A1 (n_1585), .B0 (n_1901), .C0
       (n_5333), .Y (n_5425));
  OAI211X1 g174966__6260(.A0 (\genblk2.pcpi_div_minus_2470_59_n_487 ),
       .A1 (n_1585), .B0 (n_1900), .C0 (n_5332), .Y (n_5424));
  OAI211X1 g174967__4319(.A0 (n_725), .A1 (n_1585), .B0 (n_1899), .C0
       (n_5331), .Y (n_5423));
  OAI211X1 g174968__8428(.A0 (\genblk2.pcpi_div_minus_2470_59_n_477 ),
       .A1 (n_1585), .B0 (n_1898), .C0 (n_5330), .Y (n_5422));
  OAI211X1 g174969__5526(.A0 (n_756), .A1 (n_1585), .B0 (n_1897), .C0
       (n_5329), .Y (n_5421));
  OAI211X1 g174970__6783(.A0 (\genblk2.pcpi_div_minus_2470_59_n_474 ),
       .A1 (n_1585), .B0 (n_1896), .C0 (n_5328), .Y (n_5420));
  OAI211X1 g174971__3680(.A0 (n_746), .A1 (n_1585), .B0 (n_1895), .C0
       (n_5327), .Y (n_5419));
  OAI211X1 g174972__1617(.A0 (n_714), .A1 (n_1585), .B0 (n_1893), .C0
       (n_5325), .Y (n_5418));
  OAI211X1 g174973__2802(.A0 (\genblk2.pcpi_div_minus_2470_59_n_492 ),
       .A1 (n_1585), .B0 (n_1894), .C0 (n_5326), .Y (n_5417));
  OAI211X1 g174974__1705(.A0 (\genblk2.pcpi_div_minus_2470_59_n_502 ),
       .A1 (n_1585), .B0 (n_1892), .C0 (n_5324), .Y (n_5416));
  OAI211X1 g174975__5122(.A0 (n_751), .A1 (n_1585), .B0 (n_1891), .C0
       (n_5323), .Y (n_5415));
  OAI211X1 g174976__8246(.A0 (\genblk2.pcpi_div_minus_2470_59_n_498 ),
       .A1 (n_1585), .B0 (n_1890), .C0 (n_5322), .Y (n_5414));
  OAI211X1 g174977__7098(.A0 (n_572), .A1 (n_1585), .B0 (n_1889), .C0
       (n_5321), .Y (n_5413));
  OAI211X1 g174978__6131(.A0 (\genblk2.pcpi_div_minus_2470_59_n_499 ),
       .A1 (n_1585), .B0 (n_1888), .C0 (n_5320), .Y (n_5412));
  OAI211X1 g174979__1881(.A0 (n_635), .A1 (n_1585), .B0 (n_1887), .C0
       (n_5319), .Y (n_5411));
  OAI211X1 g174980__5115(.A0 (\genblk2.pcpi_div_minus_2470_59_n_481 ),
       .A1 (n_1585), .B0 (n_1886), .C0 (n_5318), .Y (n_5410));
  OAI211X1 g174981__7482(.A0 (n_726), .A1 (n_1585), .B0 (n_1884), .C0
       (n_5317), .Y (n_5409));
  OAI211X1 g174982__4733(.A0 (\genblk2.pcpi_div_minus_2470_59_n_485 ),
       .A1 (n_1585), .B0 (n_1883), .C0 (n_5316), .Y (n_5408));
  OAI211X1 g174983__6161(.A0 (\genblk2.pcpi_div_minus_2470_59_n_500 ),
       .A1 (n_1585), .B0 (n_1882), .C0 (n_5314), .Y (n_5407));
  OAI211X1 g174984__9315(.A0 (\genblk2.pcpi_div_minus_2470_59_n_483 ),
       .A1 (n_1585), .B0 (n_1881), .C0 (n_5310), .Y (n_5406));
  OAI211X1 g174985__9945(.A0 (n_722), .A1 (n_1585), .B0 (n_1880), .C0
       (n_5309), .Y (n_5405));
  OAI211X1 g174986__2883(.A0 (\genblk2.pcpi_div_minus_2470_59_n_488 ),
       .A1 (n_1585), .B0 (n_1879), .C0 (n_5308), .Y (n_5404));
  OAI211X1 g174987__2346(.A0 (n_760), .A1 (n_1585), .B0 (n_5307), .C0
       (n_1878), .Y (n_5403));
  OAI211X1 g174988__1666(.A0 (\genblk2.pcpi_div_minus_2470_59_n_479 ),
       .A1 (n_1585), .B0 (n_5306), .C0 (n_1877), .Y (n_5402));
  OAI211X1 g174989__7410(.A0 (n_721), .A1 (n_1585), .B0 (n_5305), .C0
       (n_1876), .Y (n_5401));
  NAND2X1 g174990__6417(.A (n_2109), .B (n_5315), .Y (n_5400));
  OAI2BB1X1 g174991__5477(.A0N (\genblk2.pcpi_div_divisor [31]), .A1N
       (n_5266), .B0 (n_5334), .Y (n_5399));
  OAI2BB1X1 g174992__2398(.A0N (n_434), .A1N (\genblk2.pcpi_div_n_1998
       ), .B0 (n_5303), .Y (n_5398));
  AO21X2 g175024__8428(.A0 (n_1366), .A1 (n_5269), .B0 (n_444), .Y
       (n_5431));
  AO22X1 g175025__5526(.A0 (\genblk2.pcpi_div_divisor [23]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [22]), .B1 (n_5266), .Y
       (n_5366));
  AO22X1 g175026__6783(.A0 (\genblk2.pcpi_div_divisor [1]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [0]), .B1 (n_5266), .Y
       (n_5365));
  AO22X1 g175027__3680(.A0 (\genblk2.pcpi_div_divisor [2]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [1]), .B1 (n_5266), .Y
       (n_5364));
  AO22X1 g175028__1617(.A0 (\genblk2.pcpi_div_divisor [3]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [2]), .B1 (n_5266), .Y
       (n_5363));
  AO22X1 g175029__2802(.A0 (\genblk2.pcpi_div_divisor [4]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [3]), .B1 (n_5266), .Y
       (n_5362));
  AO22X1 g175030__1705(.A0 (\genblk2.pcpi_div_divisor [5]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [4]), .B1 (n_5266), .Y
       (n_5361));
  AO22X1 g175031__5122(.A0 (\genblk2.pcpi_div_divisor [6]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [5]), .B1 (n_5266), .Y
       (n_5360));
  AO22X1 g175032__8246(.A0 (\genblk2.pcpi_div_divisor [7]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [6]), .B1 (n_5266), .Y
       (n_5359));
  AO22X1 g175033__7098(.A0 (\genblk2.pcpi_div_divisor [8]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [7]), .B1 (n_5266), .Y
       (n_5358));
  AO22X1 g175034__6131(.A0 (\genblk2.pcpi_div_divisor [9]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [8]), .B1 (n_5266), .Y
       (n_5357));
  AO22X1 g175035__1881(.A0 (\genblk2.pcpi_div_divisor [10]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [9]), .B1 (n_5266), .Y
       (n_5356));
  AO22X1 g175036__5115(.A0 (\genblk2.pcpi_div_divisor [11]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [10]), .B1 (n_5266), .Y
       (n_5355));
  AO22X1 g175037__7482(.A0 (\genblk2.pcpi_div_divisor [12]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [11]), .B1 (n_5266), .Y
       (n_5354));
  AO22X1 g175038__4733(.A0 (\genblk2.pcpi_div_divisor [13]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [12]), .B1 (n_5266), .Y
       (n_5353));
  AO22X1 g175039__6161(.A0 (\genblk2.pcpi_div_divisor [14]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [13]), .B1 (n_5266), .Y
       (n_5352));
  AO22X1 g175040__9315(.A0 (\genblk2.pcpi_div_divisor [15]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [14]), .B1 (n_5266), .Y
       (n_5351));
  AO22X1 g175041__9945(.A0 (\genblk2.pcpi_div_divisor [17]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [16]), .B1 (n_5266), .Y
       (n_5350));
  AO22X1 g175042__2883(.A0 (\genblk2.pcpi_div_divisor [16]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [15]), .B1 (n_5266), .Y
       (n_5349));
  AO22X1 g175043__2346(.A0 (\genblk2.pcpi_div_divisor [18]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [17]), .B1 (n_5266), .Y
       (n_5348));
  AO22X1 g175044__1666(.A0 (\genblk2.pcpi_div_divisor [19]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [18]), .B1 (n_5266), .Y
       (n_5347));
  AO22X1 g175045__7410(.A0 (\genblk2.pcpi_div_divisor [20]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [19]), .B1 (n_5266), .Y
       (n_5346));
  AO22X1 g175046__6417(.A0 (\genblk2.pcpi_div_divisor [21]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [20]), .B1 (n_5266), .Y
       (n_5345));
  AO22X1 g175047__5477(.A0 (\genblk2.pcpi_div_divisor [22]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [21]), .B1 (n_5266), .Y
       (n_5344));
  OAI2BB1X1 g175048__2398(.A0N (\genblk2.pcpi_div_quotient_msk [31]),
       .A1N (n_5266), .B0 (n_954), .Y (n_5343));
  AO22X1 g175049__5107(.A0 (\genblk2.pcpi_div_divisor [24]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [23]), .B1 (n_5266), .Y
       (n_5342));
  AO22X1 g175050__6260(.A0 (\genblk2.pcpi_div_divisor [25]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [24]), .B1 (n_5266), .Y
       (n_5341));
  AO22X1 g175051__4319(.A0 (\genblk2.pcpi_div_divisor [26]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [25]), .B1 (n_5266), .Y
       (n_5340));
  AO22X1 g175052__8428(.A0 (\genblk2.pcpi_div_divisor [27]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [26]), .B1 (n_5266), .Y
       (n_5339));
  AO22X1 g175053__5526(.A0 (\genblk2.pcpi_div_divisor [28]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [27]), .B1 (n_5266), .Y
       (n_5338));
  AO22X1 g175054__6783(.A0 (\genblk2.pcpi_div_divisor [29]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [28]), .B1 (n_5266), .Y
       (n_5337));
  AO22X1 g175055__3680(.A0 (\genblk2.pcpi_div_divisor [30]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [29]), .B1 (n_5266), .Y
       (n_5336));
  AO22X1 g175056__1617(.A0 (\genblk2.pcpi_div_divisor [31]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [30]), .B1 (n_5266), .Y
       (n_5335));
  AOI22X1 g175057__2802(.A0 (\genblk2.pcpi_div_divisor [32]), .A1
       (n_5264), .B0 (\reg_op2[0]_9669 ), .B1 (n_668), .Y (n_5334));
  AOI22X1 g175058__1705(.A0 (\genblk2.pcpi_div_divisor [33]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [32]), .B1 (n_5266), .Y
       (n_5333));
  AOI22X1 g175059__5122(.A0 (\genblk2.pcpi_div_divisor [34]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [33]), .B1 (n_5266), .Y
       (n_5332));
  AOI22X1 g175060__8246(.A0 (\genblk2.pcpi_div_divisor [35]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [34]), .B1 (n_5266), .Y
       (n_5331));
  AOI22X1 g175061__7098(.A0 (\genblk2.pcpi_div_divisor [36]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [35]), .B1 (n_5266), .Y
       (n_5330));
  AOI22X1 g175062__6131(.A0 (\genblk2.pcpi_div_divisor [37]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [36]), .B1 (n_5266), .Y
       (n_5329));
  AOI22X1 g175063__1881(.A0 (\genblk2.pcpi_div_divisor [38]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [37]), .B1 (n_5266), .Y
       (n_5328));
  AOI22X1 g175064__5115(.A0 (\genblk2.pcpi_div_divisor [39]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [38]), .B1 (n_5266), .Y
       (n_5327));
  AOI22X1 g175065__7482(.A0 (\genblk2.pcpi_div_divisor [40]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [39]), .B1 (n_5266), .Y
       (n_5326));
  AOI22X1 g175066__4733(.A0 (\genblk2.pcpi_div_divisor [41]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [40]), .B1 (n_5266), .Y
       (n_5325));
  AOI22X1 g175067__6161(.A0 (\genblk2.pcpi_div_divisor [42]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [41]), .B1 (n_5266), .Y
       (n_5324));
  AOI22X1 g175068__9315(.A0 (\genblk2.pcpi_div_divisor [43]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [42]), .B1 (n_5266), .Y
       (n_5323));
  AOI22X1 g175069__9945(.A0 (\genblk2.pcpi_div_divisor [44]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [43]), .B1 (n_5266), .Y
       (n_5322));
  AOI22X1 g175070__2883(.A0 (\genblk2.pcpi_div_divisor [45]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [44]), .B1 (n_5266), .Y
       (n_5321));
  AOI22X1 g175071__2346(.A0 (\genblk2.pcpi_div_divisor [46]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [45]), .B1 (n_5266), .Y
       (n_5320));
  AOI22X1 g175073__1666(.A0 (\genblk2.pcpi_div_divisor [47]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [46]), .B1 (n_5266), .Y
       (n_5319));
  AOI22X1 g175074__7410(.A0 (\genblk2.pcpi_div_divisor [48]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [47]), .B1 (n_5266), .Y
       (n_5318));
  AOI22X1 g175075__6417(.A0 (\genblk2.pcpi_div_divisor [49]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [48]), .B1 (n_5266), .Y
       (n_5317));
  AOI22X1 g175076__5477(.A0 (\genblk2.pcpi_div_divisor [50]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [49]), .B1 (n_5266), .Y
       (n_5316));
  AOI22X1 g175077__2398(.A0 (\genblk2.pcpi_div_divisor [51]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [50]), .B1 (n_5266), .Y
       (n_5315));
  AOI22X1 g175078__5107(.A0 (\genblk2.pcpi_div_divisor [52]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [51]), .B1 (n_5266), .Y
       (n_5314));
  AOI22X1 g175079__6260(.A0 (\genblk2.pcpi_div_divisor [53]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [52]), .B1 (n_5266), .Y
       (n_5313));
  AOI22X1 g175080__4319(.A0 (\genblk2.pcpi_div_divisor [54]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [53]), .B1 (n_5266), .Y
       (n_5312));
  AOI22X1 g175081__8428(.A0 (\genblk2.pcpi_div_divisor [55]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [54]), .B1 (n_5266), .Y
       (n_5311));
  AOI22X1 g175082__5526(.A0 (\genblk2.pcpi_div_divisor [56]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [55]), .B1 (n_5266), .Y
       (n_5310));
  AOI22X1 g175083__6783(.A0 (\genblk2.pcpi_div_divisor [57]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [56]), .B1 (n_5266), .Y
       (n_5309));
  AOI22X1 g175084__3680(.A0 (\genblk2.pcpi_div_divisor [58]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [57]), .B1 (n_5266), .Y
       (n_5308));
  AOI22X1 g175085__1617(.A0 (\genblk2.pcpi_div_divisor [59]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [58]), .B1 (n_5266), .Y
       (n_5307));
  AOI22X1 g175086__2802(.A0 (\genblk2.pcpi_div_divisor [60]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [59]), .B1 (n_5266), .Y
       (n_5306));
  AOI22X1 g175087__1705(.A0 (\genblk2.pcpi_div_divisor [61]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [60]), .B1 (n_5266), .Y
       (n_5305));
  AOI22X1 g175088__5122(.A0 (\genblk2.pcpi_div_divisor [62]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_divisor [61]), .B1 (n_5266), .Y
       (n_5304));
  AOI22X1 g175089__8246(.A0 (\genblk2.pcpi_div_divisor [62]), .A1
       (n_5266), .B0 (\reg_op2[31]_9700 ), .B1 (n_1584), .Y (n_5303));
  AO22X1 g175090__7098(.A0 (\genblk2.pcpi_div_quotient_msk [1]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_quotient_msk [0]), .B1
       (n_5266), .Y (n_5302));
  AO22X1 g175091__6131(.A0 (\genblk2.pcpi_div_quotient_msk [2]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_quotient_msk [1]), .B1
       (n_5266), .Y (n_5301));
  AO22X1 g175092__1881(.A0 (\genblk2.pcpi_div_quotient_msk [3]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_quotient_msk [2]), .B1
       (n_5266), .Y (n_5300));
  AO22X1 g175093__5115(.A0 (\genblk2.pcpi_div_quotient_msk [4]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_quotient_msk [3]), .B1
       (n_5266), .Y (n_5299));
  AO22X1 g175094__7482(.A0 (\genblk2.pcpi_div_quotient_msk [5]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_quotient_msk [4]), .B1
       (n_5266), .Y (n_5298));
  AO22X1 g175095__4733(.A0 (\genblk2.pcpi_div_quotient_msk [8]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_quotient_msk [7]), .B1
       (n_5266), .Y (n_5297));
  AO22X1 g175096__6161(.A0 (\genblk2.pcpi_div_quotient_msk [9]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_quotient_msk [8]), .B1
       (n_5266), .Y (n_5296));
  AO22X1 g175097__9315(.A0 (\genblk2.pcpi_div_quotient_msk [7]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_quotient_msk [6]), .B1
       (n_5266), .Y (n_5295));
  AO22X1 g175098__9945(.A0 (\genblk2.pcpi_div_quotient_msk [10]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_quotient_msk [9]), .B1
       (n_5266), .Y (n_5294));
  AO22X1 g175099__2883(.A0 (\genblk2.pcpi_div_quotient_msk [11]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_quotient_msk [10]), .B1
       (n_5266), .Y (n_5293));
  AO22X1 g175100__2346(.A0 (\genblk2.pcpi_div_quotient_msk [12]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_quotient_msk [11]), .B1
       (n_5266), .Y (n_5292));
  AO22X1 g175101__1666(.A0 (\genblk2.pcpi_div_quotient_msk [6]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_quotient_msk [5]), .B1
       (n_5266), .Y (n_5291));
  AO22X1 g175102__7410(.A0 (\genblk2.pcpi_div_quotient_msk [13]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_quotient_msk [12]), .B1
       (n_5266), .Y (n_5290));
  AO22X1 g175103__6417(.A0 (\genblk2.pcpi_div_quotient_msk [14]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_quotient_msk [13]), .B1
       (n_5266), .Y (n_5289));
  AO22X1 g175104__5477(.A0 (\genblk2.pcpi_div_quotient_msk [15]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_quotient_msk [14]), .B1
       (n_5266), .Y (n_5288));
  AO22X1 g175105__2398(.A0 (\genblk2.pcpi_div_quotient_msk [16]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_quotient_msk [15]), .B1
       (n_5266), .Y (n_5287));
  AO22X1 g175106__5107(.A0 (\genblk2.pcpi_div_quotient_msk [17]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_quotient_msk [16]), .B1
       (n_5266), .Y (n_5286));
  AO22X1 g175107__6260(.A0 (\genblk2.pcpi_div_quotient_msk [18]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_quotient_msk [17]), .B1
       (n_5266), .Y (n_5285));
  AO22X1 g175108__4319(.A0 (\genblk2.pcpi_div_quotient_msk [19]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_quotient_msk [18]), .B1
       (n_5266), .Y (n_5284));
  AO22X1 g175109__8428(.A0 (\genblk2.pcpi_div_quotient_msk [20]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_quotient_msk [19]), .B1
       (n_5266), .Y (n_5283));
  AO22X1 g175110__5526(.A0 (\genblk2.pcpi_div_quotient_msk [21]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_quotient_msk [20]), .B1
       (n_5266), .Y (n_5282));
  AO22X1 g175111__6783(.A0 (\genblk2.pcpi_div_quotient_msk [23]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_quotient_msk [22]), .B1
       (n_5266), .Y (n_5281));
  AO22X1 g175112__3680(.A0 (\genblk2.pcpi_div_quotient_msk [24]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_quotient_msk [23]), .B1
       (n_5266), .Y (n_5280));
  AO22X1 g175113__1617(.A0 (\genblk2.pcpi_div_quotient_msk [22]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_quotient_msk [21]), .B1
       (n_5266), .Y (n_5279));
  AO22X1 g175114__2802(.A0 (\genblk2.pcpi_div_quotient_msk [25]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_quotient_msk [24]), .B1
       (n_5266), .Y (n_5278));
  AO22X1 g175115__1705(.A0 (\genblk2.pcpi_div_quotient_msk [26]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_quotient_msk [25]), .B1
       (n_5266), .Y (n_5277));
  AO22X1 g175116__5122(.A0 (\genblk2.pcpi_div_quotient_msk [27]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_quotient_msk [26]), .B1
       (n_5266), .Y (n_5276));
  AO22X1 g175117__8246(.A0 (\genblk2.pcpi_div_quotient_msk [28]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_quotient_msk [27]), .B1
       (n_5266), .Y (n_5275));
  AO22X1 g175118__7098(.A0 (\genblk2.pcpi_div_quotient_msk [29]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_quotient_msk [28]), .B1
       (n_5266), .Y (n_5274));
  AO22X1 g175119__6131(.A0 (\genblk2.pcpi_div_quotient_msk [30]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_quotient_msk [29]), .B1
       (n_5266), .Y (n_5273));
  AO22X1 g175120__1881(.A0 (\genblk2.pcpi_div_quotient_msk [31]), .A1
       (n_5264), .B0 (\genblk2.pcpi_div_quotient_msk [30]), .B1
       (n_5266), .Y (n_5272));
  AND2X2 g175122__5115(.A (\genblk2.pcpi_div_n_314 ), .B (n_5264), .Y
       (n_444));
  INVX2 g175123(.A (n_5269), .Y (n_5270));
  OAI21X1 g175124__7482(.A0 (n_544), .A1 (n_1365), .B0 (n_5263), .Y
       (n_5268));
  AOI221X1 g175125__4733(.A0 (n_2297), .A1 (n_5257), .B0
       (\reg_op2[24]_9693 ), .B1 (n_713), .C0 (n_876), .Y (n_5267));
  AOI21X1 g175126__6161(.A0 (\genblk2.pcpi_div_n_4742 ), .A1 (n_609),
       .B0 (n_5266), .Y (n_5269));
  NOR2X1 g175127__9315(.A (n_544), .B (n_5260), .Y (n_5265));
  OR2X4 g175128__9945(.A (n_544), .B (n_5261), .Y (n_5266));
  NAND3BXL g175129__2883(.AN (n_294), .B (\genblk2.pcpi_div_running ),
       .C (n_1365), .Y (n_5263));
  OAI2BB1X1 g175130__2346(.A0N (\genblk2.pcpi_div_instr_rem ), .A1N
       (\reg_op1[31]_9668 ), .B0 (n_5259), .Y (n_5262));
  AND3X4 g175131__1666(.A (\genblk2.pcpi_div_n_4742 ), .B (n_543), .C
       (n_706), .Y (n_5264));
  INVX1 g175133(.A (n_5260), .Y (n_5261));
  OAI211X1 g175134__7410(.A0 (\reg_op2[31]_9700 ), .A1 (n_5236), .B0
       (\genblk2.pcpi_div_instr_div ), .C0 (n_11691), .Y (n_5259));
  NAND2X1 g175135__6417(.A (\genblk2.pcpi_div_n_4742 ), .B (n_294), .Y
       (n_5260));
  AOI221X1 g175146__5477(.A0 (n_138), .A1 (n_812), .B0 (n_154), .B1
       (n_5239), .C0 (n_1921), .Y (n_5257));
  MX2X1 g175147__2398(.A (\reg_op1[29]_9666 ), .B (n_5240), .S0
       (n_321), .Y (n_5256));
  NOR4X1 g175148__5107(.A (\genblk2.pcpi_div_quotient_msk [31]), .B
       (\genblk2.pcpi_div_quotient_msk [25]), .C
       (\genblk2.pcpi_div_quotient_msk [17]), .D (n_5227), .Y (n_294));
  MX2X1 g175155__6260(.A (\reg_op1[4]_9641 ), .B (n_5226), .S0
       (n_2489), .Y (n_5255));
  MX2X1 g175156__4319(.A (\reg_op1[9]_9646 ), .B (n_5223), .S0
       (n_2489), .Y (n_5254));
  MX2X1 g175157__8428(.A (\reg_op1[8]_9645 ), .B (n_5224), .S0 (n_321),
       .Y (n_5253));
  MX2X1 g175158__5526(.A (\reg_op1[5]_9642 ), .B (n_5225), .S0
       (n_2489), .Y (n_5252));
  MX2X1 g175166__6783(.A (\reg_op1[24]_9661 ), .B (n_5218), .S0
       (n_321), .Y (n_5251));
  MX2X1 g175167__3680(.A (\reg_op1[11]_9648 ), .B (n_5222), .S0
       (n_2489), .Y (n_5250));
  MX2X1 g175168__1617(.A (\reg_op1[12]_9649 ), .B (n_5220), .S0
       (n_321), .Y (n_5249));
  MX2X1 g175169__2802(.A (\reg_op1[13]_9650 ), .B (n_5219), .S0
       (n_2489), .Y (n_5248));
  MX2X1 g175170__1705(.A (\reg_op1[17]_9654 ), .B (n_5217), .S0
       (n_321), .Y (n_5247));
  MX2X1 g175171__5122(.A (\reg_op1[10]_9647 ), .B (n_5230), .S0
       (n_2489), .Y (n_5246));
  MX2X1 g175172__8246(.A (\reg_op1[26]_9663 ), .B (n_5216), .S0
       (n_321), .Y (n_5245));
  MX2X1 g175173__7098(.A (\reg_op1[27]_9664 ), .B (n_5221), .S0
       (n_321), .Y (n_5244));
  OAI22X1 g175174__6131(.A0 (n_5215), .A1 (n_693), .B0 (n_744), .B1
       (n_2489), .Y (n_5243));
  MX2X1 g175175__1881(.A (\reg_op1[28]_9665 ), .B (n_5228), .S0
       (n_2489), .Y (n_5242));
  MX2X1 g175176__5115(.A (\reg_op1[23]_9660 ), .B (n_5213), .S0
       (n_321), .Y (n_5241));
  NAND4XL g175177__7482(.A (n_1640), .B (n_2197), .C (n_5181), .D
       (n_2196), .Y (n_5240));
  NOR4X1 g175178__4733(.A (n_825), .B (n_1358), .C (n_1635), .D
       (n_5194), .Y (n_5239));
  MX2X1 g175179__6161(.A (n_5203), .B (\reg_op1[15]_9652 ), .S0
       (n_693), .Y (n_5238));
  MX2X1 g175180(.A (n_5212), .B (\reg_op1[6]_9643 ), .S0 (n_693), .Y
       (n_5237));
  NAND4XL g175183(.A (\genblk2.pcpi_div_minus_2470_59_n_485 ), .B
       (\genblk2.pcpi_div_minus_2470_59_n_481 ), .C
       (\genblk2.pcpi_div_minus_2470_59_n_479 ), .D (n_5193), .Y
       (n_5236));
  NAND4XL g175184(.A (n_2424), .B (n_2606), .C (n_5081), .D (n_5177),
       .Y (n_5235));
  MX2X1 g175185(.A (n_5210), .B (reg_op1[0]), .S0 (n_693), .Y (n_5234));
  OAI22X1 g175186(.A0 (n_693), .A1 (n_5208), .B0 (n_747), .B1 (n_321),
       .Y (n_5233));
  OAI22X1 g175187(.A0 (n_693), .A1 (n_5207), .B0 (n_576), .B1 (n_2489),
       .Y (n_5232));
  OAI22X1 g175188(.A0 (n_5209), .A1 (n_693), .B0 (n_565), .B1 (n_321),
       .Y (n_5231));
  NAND3X1 g175189(.A (n_2209), .B (n_2355), .C (n_5190), .Y (n_5230));
  NAND2X1 g175190(.A (n_5114), .B (n_5205), .Y (n_5229));
  NAND4XL g175191(.A (n_1640), .B (n_2158), .C (n_5182), .D (n_2367),
       .Y (n_5228));
  OR4X1 g175192(.A (\genblk2.pcpi_div_quotient_msk [18]), .B
       (\genblk2.pcpi_div_quotient_msk [19]), .C
       (\genblk2.pcpi_div_quotient_msk [20]), .D (n_5172), .Y (n_5227));
  NAND3X1 g175193(.A (n_2216), .B (n_2386), .C (n_5192), .Y (n_5226));
  NAND3X1 g175194(.A (n_2214), .B (n_2365), .C (n_5191), .Y (n_5225));
  NAND3X1 g175195(.A (n_2211), .B (n_2357), .C (n_5201), .Y (n_5224));
  NAND3X1 g175196(.A (n_2210), .B (n_2356), .C (n_5202), .Y (n_5223));
  NAND3X1 g175199(.A (n_2208), .B (n_2359), .C (n_5189), .Y (n_5222));
  NAND3X1 g175200(.A (n_2215), .B (n_5183), .C (n_2368), .Y (n_5221));
  NAND3X1 g175201(.A (n_2207), .B (n_2358), .C (n_5188), .Y (n_5220));
  NAND3X1 g175202(.A (n_2206), .B (n_2360), .C (n_5187), .Y (n_5219));
  NAND3X1 g175203(.A (n_2200), .B (n_5185), .C (n_2370), .Y (n_5218));
  NAND3X1 g175204(.A (n_2202), .B (n_5186), .C (n_2361), .Y (n_5217));
  NAND3X1 g175205(.A (n_2212), .B (n_5184), .C (n_2369), .Y (n_5216));
  AOI221X1 g175206(.A0 (\reg_op1[8]_9645 ), .A1 (n_550), .B0
       (\reg_op1[11]_9648 ), .B1 (n_332), .C0 (n_5211), .Y (n_5215));
  OAI22X1 g175207(.A0 (n_693), .A1 (n_5195), .B0 (n_625), .B1 (n_2489),
       .Y (n_5214));
  OAI211X1 g175208(.A0 (n_576), .A1 (n_1940), .B0 (n_2177), .C0
       (n_5199), .Y (n_5213));
  NAND3X1 g175209(.A (n_2213), .B (n_2364), .C (n_5164), .Y (n_5212));
  NAND4XL g175218(.A (n_2159), .B (n_4750), .C (n_4749), .D (n_5165),
       .Y (n_5211));
  OAI211X1 g175219(.A0 (n_565), .A1 (n_677), .B0 (n_2205), .C0
       (n_5171), .Y (n_5210));
  AOI221X1 g175220(.A0 (n_1932), .A1 (n_5132), .B0 (\reg_op1[5]_9642 ),
       .B1 (n_332), .C0 (n_2180), .Y (n_5209));
  AOI221X1 g175221(.A0 (\reg_op1[20]_9657 ), .A1 (n_550), .B0
       (\reg_op1[23]_9660 ), .B1 (n_332), .C0 (n_5197), .Y (n_5208));
  AOI221X1 g175222(.A0 (\reg_op1[23]_9660 ), .A1 (n_550), .B0
       (\reg_op1[26]_9663 ), .B1 (n_332), .C0 (n_5196), .Y (n_5207));
  OAI22X1 g175223(.A0 (n_693), .A1 (n_5166), .B0 (n_634), .B1 (n_321),
       .Y (n_5206));
  AOI221X1 g175224(.A0 (n_317), .A1 (n_5134), .B0 (mem_rdata_q[25]),
       .B1 (n_5025), .C0 (n_5106), .Y (n_5205));
  OAI22X1 g175225(.A0 (n_693), .A1 (n_5173), .B0 (n_637), .B1 (n_321),
       .Y (n_5204));
  NAND3X1 g175226(.A (n_2204), .B (n_2362), .C (n_5163), .Y (n_5203));
  AOI22X1 g175227(.A0 (cpu_state[5]), .A1 (n_5141), .B0
       (\reg_op1[13]_9650 ), .B1 (n_332), .Y (n_5202));
  AOI22X1 g175228(.A0 (cpu_state[5]), .A1 (n_5142), .B0
       (\reg_op1[12]_9649 ), .B1 (n_332), .Y (n_5201));
  OAI211X1 g175229(.A0 (n_1806), .A1 (n_301), .B0 (n_5115), .C0
       (n_5136), .Y (n_5200));
  AOI221X1 g175230(.A0 (\cpuregs[5] [23]), .A1 (n_11748), .B0 (n_833),
       .B1 (n_6937), .C0 (n_5159), .Y (n_5199));
  NAND4XL g175231(.A (n_2535), .B (n_5114), .C (n_5065), .D (n_5102),
       .Y (n_5198));
  OAI211X1 g175232(.A0 (n_625), .A1 (n_1940), .B0 (n_5152), .C0
       (n_4857), .Y (n_5197));
  OAI211X1 g175233(.A0 (n_637), .A1 (n_1940), .B0 (n_5158), .C0
       (n_4856), .Y (n_5196));
  AOI221X1 g175234(.A0 (\reg_op1[19]_9656 ), .A1 (n_550), .B0
       (\reg_op1[22]_9659 ), .B1 (n_332), .C0 (n_5167), .Y (n_5195));
  AOI32X1 g175235(.A0 (n_862), .A1 (n_855), .A2 (n_5146), .B0 (n_855),
       .B1 (n_1308), .Y (n_5194));
  NOR4X1 g175236(.A (\reg_op2[19]_9688 ), .B (\reg_op2[17]_9686 ), .C
       (\reg_op2[1]_9670 ), .D (n_5107), .Y (n_5193));
  AOI22X1 g175237(.A0 (cpu_state[5]), .A1 (n_5143), .B0
       (\reg_op1[8]_9645 ), .B1 (n_332), .Y (n_5192));
  AOI22X1 g175238(.A0 (cpu_state[5]), .A1 (n_5131), .B0
       (\reg_op1[9]_9646 ), .B1 (n_332), .Y (n_5191));
  AOI22X1 g175244(.A0 (cpu_state[5]), .A1 (n_5130), .B0
       (\reg_op1[14]_9651 ), .B1 (n_332), .Y (n_5190));
  AOI22X1 g175245(.A0 (cpu_state[5]), .A1 (n_5140), .B0
       (\reg_op1[15]_9652 ), .B1 (n_332), .Y (n_5189));
  AOI22X1 g175246(.A0 (cpu_state[5]), .A1 (n_5139), .B0
       (\reg_op1[16]_9653 ), .B1 (n_332), .Y (n_5188));
  AOI22X1 g175247(.A0 (cpu_state[5]), .A1 (n_5129), .B0
       (\reg_op1[17]_9654 ), .B1 (n_332), .Y (n_5187));
  AOI22X1 g175248(.A0 (cpu_state[5]), .A1 (n_5138), .B0
       (\reg_op1[21]_9658 ), .B1 (n_332), .Y (n_5186));
  AOI22X1 g175249(.A0 (cpu_state[5]), .A1 (n_5137), .B0
       (\reg_op1[28]_9665 ), .B1 (n_332), .Y (n_5185));
  AOI22X1 g175250(.A0 (cpu_state[5]), .A1 (n_5128), .B0
       (\reg_op1[30]_9667 ), .B1 (n_332), .Y (n_5184));
  AOI22X1 g175251(.A0 (cpu_state[5]), .A1 (n_5127), .B0
       (\reg_op1[31]_9668 ), .B1 (n_332), .Y (n_5183));
  AOI22X1 g175252(.A0 (cpu_state[5]), .A1 (n_5126), .B0 (reg_pc[28]),
       .B1 (n_547), .Y (n_5182));
  AOI22X1 g175253(.A0 (cpu_state[5]), .A1 (n_5145), .B0
       (\reg_op1[30]_9667 ), .B1 (n_550), .Y (n_5181));
  OAI22X1 g175254(.A0 (n_693), .A1 (n_5153), .B0 (n_627), .B1 (n_2489),
       .Y (n_5180));
  OAI22X1 g175255(.A0 (n_693), .A1 (n_5154), .B0 (n_718), .B1 (n_321),
       .Y (n_5179));
  OAI221X1 g175256(.A0 (n_2131), .A1 (n_301), .B0 (n_680), .B1 (n_308),
       .C0 (n_5162), .Y (n_5178));
  AOI221X1 g175257(.A0 (n_2137), .A1 (n_5116), .B0 (n_439), .B1
       (n_5119), .C0 (n_5093), .Y (n_5177));
  MX2X1 g175258(.A (n_5150), .B (\reg_op1[14]_9651 ), .S0 (n_693), .Y
       (n_5176));
  MX2X1 g175259(.A (n_5148), .B (\reg_op1[16]_9653 ), .S0 (n_693), .Y
       (n_5175));
  MX2X1 g175260(.A (n_5147), .B (\reg_op1[25]_9662 ), .S0 (n_693), .Y
       (n_5174));
  AOI221X1 g175261(.A0 (\reg_op1[25]_9662 ), .A1 (n_332), .B0
       (\reg_op1[17]_9654 ), .B1 (n_1944), .C0 (n_5155), .Y (n_5173));
  OR4X1 g175262(.A (\genblk2.pcpi_div_quotient_msk [21]), .B
       (\genblk2.pcpi_div_quotient_msk [22]), .C
       (\genblk2.pcpi_div_quotient_msk [1]), .D (n_5092), .Y (n_5172));
  NAND2X1 g175263(.A (cpu_state[5]), .B (n_5133), .Y (n_5171));
  NAND2X1 g175264(.A (n_5114), .B (n_5157), .Y (n_5170));
  NAND2X1 g175265(.A (n_5114), .B (n_5156), .Y (n_5169));
  NAND2X1 g175266(.A (n_5115), .B (n_5135), .Y (n_5168));
  OAI222X1 g175270(.A0 (n_715), .A1 (n_1940), .B0 (n_1935), .B1
       (n_5086), .C0 (n_624), .C1 (n_1943), .Y (n_5167));
  AOI211XL g175271(.A0 (n_833), .A1 (n_6940), .B0 (n_2389), .C0
       (n_5124), .Y (n_5166));
  AOI222X1 g175272(.A0 (n_833), .A1 (n_6953), .B0 (cpu_state[5]), .B1
       (n_5088), .C0 (reg_pc[7]), .C1 (n_547), .Y (n_5165));
  AOI22X1 g175273(.A0 (cpu_state[5]), .A1 (n_5100), .B0
       (\reg_op1[10]_9647 ), .B1 (n_332), .Y (n_5164));
  AOI22X1 g175274(.A0 (cpu_state[5]), .A1 (n_5101), .B0
       (\reg_op1[19]_9656 ), .B1 (n_332), .Y (n_5163));
  AOI221X1 g175275(.A0 (mem_rdata_q[12]), .A1 (n_5025), .B0 (n_439),
       .B1 (n_2436), .C0 (n_5144), .Y (n_5162));
  OAI22X1 g175276(.A0 (n_5112), .A1 (n_693), .B0 (n_578), .B1 (n_321),
       .Y (n_5161));
  OAI22X1 g175277(.A0 (n_5111), .A1 (n_693), .B0 (n_577), .B1 (n_2489),
       .Y (n_5160));
  OAI211X1 g175278(.A0 (n_548), .A1 (n_5068), .B0 (n_1531), .C0
       (n_4742), .Y (n_5159));
  AOI221X1 g175279(.A0 (cpu_state[5]), .A1 (n_5055), .B0 (reg_pc[22]),
       .B1 (n_547), .C0 (n_4743), .Y (n_5158));
  AOI221X1 g175280(.A0 (n_326), .A1 (n_2585), .B0 (n_504), .B1 (n_17),
       .C0 (n_5105), .Y (n_5157));
  AOI221X1 g175281(.A0 (n_2146), .A1 (n_2585), .B0 (n_2137), .B1
       (n_2436), .C0 (n_5104), .Y (n_5156));
  OAI211X1 g175282(.A0 (n_634), .A1 (n_1940), .B0 (n_2201), .C0
       (n_5083), .Y (n_5155));
  NOR4X1 g175283(.A (n_1340), .B (n_4), .C (n_2273), .D (n_5048), .Y
       (n_5154));
  NOR2BX1 g175284(.AN (n_5110), .B (n_1340), .Y (n_5153));
  AOI221X1 g175285(.A0 (cpu_state[5]), .A1 (n_5056), .B0 (reg_pc[19]),
       .B1 (n_547), .C0 (n_4746), .Y (n_5152));
  OAI211X1 g175286(.A0 (n_1809), .A1 (n_301), .B0 (n_5052), .C0
       (n_5115), .Y (n_5151));
  OAI221X1 g175287(.A0 (n_619), .A1 (n_677), .B0 (n_625), .B1 (n_678),
       .C0 (n_5109), .Y (n_5150));
  OAI211X1 g175288(.A0 (n_984), .A1 (n_975), .B0 (n_4534), .C0
       (n_5108), .Y (n_5149));
  NAND4XL g175289(.A (n_2181), .B (n_4748), .C (n_5077), .D (n_2203),
       .Y (n_5148));
  NAND4XL g175290(.A (n_2188), .B (n_4741), .C (n_5074), .D (n_2199),
       .Y (n_5147));
  OAI2BB1X1 g175291(.A0N (n_11740), .A1N (n_5085), .B0 (n_865), .Y
       (n_5146));
  NAND4XL g175299(.A (n_4670), .B (n_4669), .C (n_4770), .D (n_5070),
       .Y (n_5145));
  OAI22X1 g175300(.A0 (n_2517), .A1 (n_5098), .B0 (n_2438), .B1
       (n_5060), .Y (n_5144));
  NAND4XL g175301(.A (n_4469), .B (n_4470), .C (n_4468), .D (n_5094),
       .Y (n_5143));
  NAND4XL g175302(.A (n_4421), .B (n_4422), .C (n_4420), .D (n_5096),
       .Y (n_5142));
  NAND4XL g175303(.A (n_4407), .B (n_4408), .C (n_4406), .D (n_5097),
       .Y (n_5141));
  NAND4XL g175304(.A (n_4382), .B (n_4383), .C (n_4381), .D (n_5080),
       .Y (n_5140));
  NAND4XL g175305(.A (n_4368), .B (n_4369), .C (n_4367), .D (n_5079),
       .Y (n_5139));
  NAND4XL g175306(.A (n_4301), .B (n_4302), .C (n_4300), .D (n_5076),
       .Y (n_5138));
  NAND4XL g175307(.A (n_4608), .B (n_4607), .C (n_4609), .D (n_5075),
       .Y (n_5137));
  AOI22X1 g175308(.A0 (n_2568), .A1 (n_5099), .B0 (mem_rdata_q[30]),
       .B1 (n_5025), .Y (n_5136));
  AOI222X1 g175309(.A0 (mem_rdata_q[29]), .A1 (n_5025), .B0 (n_1805),
       .B1 (n_705), .C0 (n_503), .C1 (n_14), .Y (n_5135));
  OAI211X1 g175310(.A0 (n_2319), .A1 (n_5060), .B0 (n_2422), .C0
       (n_2424), .Y (n_5134));
  NAND4XL g175311(.A (n_4523), .B (n_4522), .C (n_4787), .D (n_5090),
       .Y (n_5133));
  NAND4XL g175312(.A (n_4511), .B (n_4510), .C (n_4512), .D (n_5089),
       .Y (n_5132));
  NAND4XL g175313(.A (n_4456), .B (n_4455), .C (n_4784), .D (n_5095),
       .Y (n_5131));
  NAND4XL g175314(.A (n_4394), .B (n_4393), .C (n_4781), .D (n_5061),
       .Y (n_5130));
  NAND4XL g175315(.A (n_4354), .B (n_4355), .C (n_4780), .D (n_5078),
       .Y (n_5129));
  NAND4XL g175316(.A (n_4635), .B (n_4636), .C (n_4794), .D (n_5073),
       .Y (n_5128));
  NAND4XL g175317(.A (n_4646), .B (n_4647), .C (n_4772), .D (n_5072),
       .Y (n_5127));
  NAND4XL g175318(.A (n_4658), .B (n_4657), .C (n_4771), .D (n_5071),
       .Y (n_5126));
  OAI211X1 g175319(.A0 (n_679), .A1 (n_308), .B0 (n_5053), .C0
       (n_5113), .Y (n_5125));
  OAI2BB1X1 g175320(.A0N (reg_pc[20]), .A1N (n_547), .B0 (n_5087), .Y
       (n_5124));
  NAND2X1 g175321(.A (n_329), .B (n_5062), .Y (n_5123));
  NAND2X1 g175322(.A (n_329), .B (n_5063), .Y (n_5122));
  OAI211X1 g175323(.A0 (n_1954), .A1 (n_5027), .B0 (n_543), .C0
       (n_5041), .Y (n_5121));
  OAI211X1 g175324(.A0 (n_644), .A1 (n_341), .B0 (n_329), .C0 (n_5036),
       .Y (n_5120));
  OAI2BB1X1 g175325(.A0N (n_2321), .A1N (n_5059), .B0 (n_3469), .Y
       (n_5119));
  OAI211X1 g175326(.A0 (n_588), .A1 (n_341), .B0 (n_329), .C0 (n_5035),
       .Y (n_5118));
  NAND4XL g175327(.A (n_329), .B (n_3415), .C (n_4953), .D (n_5023), .Y
       (n_5117));
  NOR2X1 g175328(.A (n_325), .B (n_5098), .Y (n_5116));
  AOI32X1 g175336(.A0 (n_15), .A1 (n_3006), .A2 (n_5059), .B0 (n_438),
       .B1 (n_705), .Y (n_5113));
  AOI221X1 g175337(.A0 (n_1934), .A1 (n_5018), .B0 (\reg_op1[7]_9644 ),
       .B1 (n_332), .C0 (n_2187), .Y (n_5112));
  AOI221X1 g175338(.A0 (n_1933), .A1 (n_5019), .B0 (\reg_op1[6]_9643 ),
       .B1 (n_332), .C0 (n_2178), .Y (n_5111));
  AOI222X1 g175339(.A0 (\reg_op1[30]_9667 ), .A1 (n_1941), .B0
       (n_1930), .B1 (n_5017), .C0 (\reg_op1[27]_9664 ), .C1 (n_1944),
       .Y (n_5110));
  AOI222X1 g175340(.A0 (\reg_op1[13]_9650 ), .A1 (n_1941), .B0
       (n_1931), .B1 (n_5015), .C0 (\reg_op1[10]_9647 ), .C1 (n_1944),
       .Y (n_5109));
  AOI32X1 g175341(.A0 (n_645), .A1 (n_1339), .A2 (n_5028), .B0
       (cpu_state[7]), .B1 (n_348), .Y (n_5108));
  NAND4XL g175342(.A (n_721), .B (\genblk2.pcpi_div_minus_2470_59_n_483
       ), .C (n_760), .D (n_5013), .Y (n_5107));
  OAI22X1 g175343(.A0 (n_1804), .A1 (n_301), .B0 (n_680), .B1 (n_3249),
       .Y (n_5106));
  OAI222X1 g175344(.A0 (n_591), .A1 (n_5026), .B0 (n_1816), .B1
       (n_301), .C0 (n_686), .C1 (n_3419), .Y (n_5105));
  OAI222X1 g175345(.A0 (n_642), .A1 (n_5026), .B0 (n_1808), .B1
       (n_301), .C0 (n_682), .C1 (n_3174), .Y (n_5104));
  OAI22X1 g175346(.A0 (n_537), .A1 (n_5042), .B0 (n_558), .B1 (n_538),
       .Y (n_5103));
  AOI22X1 g175347(.A0 (n_1814), .A1 (n_705), .B0 (n_334), .B1 (n_3066),
       .Y (n_5102));
  NAND4XL g175348(.A (n_4329), .B (n_4328), .C (n_4778), .D (n_5039),
       .Y (n_5101));
  NAND4XL g175349(.A (n_4444), .B (n_4445), .C (n_4783), .D (n_5040),
       .Y (n_5100));
  OAI211X1 g175350(.A0 (n_438), .A1 (n_2599), .B0 (n_317), .C0
       (n_5059), .Y (n_5115));
  OAI211X1 g175351(.A0 (n_2997), .A1 (n_2599), .B0 (n_317), .C0
       (n_5059), .Y (n_5114));
  INVX1 g175352(.A (n_5098), .Y (n_5099));
  AOI211XL g175353(.A0 (\cpuregs[5] [9]), .A1 (n_291), .B0 (n_4795),
       .C0 (n_5007), .Y (n_5097));
  AOI211XL g175354(.A0 (\cpuregs[5] [8]), .A1 (n_291), .B0 (n_4874),
       .C0 (n_5008), .Y (n_5096));
  AOI221X1 g175355(.A0 (\cpuregs[1] [5]), .A1 (n_456), .B0
       (\cpuregs[2] [5]), .B1 (n_425), .C0 (n_5049), .Y (n_5095));
  AOI211XL g175356(.A0 (\cpuregs[5] [4]), .A1 (n_291), .B0 (n_4867),
       .C0 (n_5010), .Y (n_5094));
  NOR2X1 g175357(.A (n_2332), .B (n_5060), .Y (n_5093));
  OR4X1 g175358(.A (\genblk2.pcpi_div_quotient_msk [2]), .B
       (\genblk2.pcpi_div_quotient_msk [3]), .C
       (\genblk2.pcpi_div_quotient_msk [4]), .D (n_4986), .Y (n_5092));
  NAND2X1 g175359(.A (n_3467), .B (n_5034), .Y (n_5091));
  AOI221X1 g175360(.A0 (\cpuregs[1] [0]), .A1 (n_456), .B0
       (\cpuregs[2] [0]), .B1 (n_425), .C0 (n_5047), .Y (n_5090));
  AOI221X1 g175361(.A0 (\cpuregs[30] [1]), .A1 (n_500), .B0
       (\cpuregs[31] [1]), .B1 (n_476), .C0 (n_5057), .Y (n_5089));
  NAND4XL g175362(.A (n_4114), .B (n_4782), .C (n_4912), .D (n_4983),
       .Y (n_5088));
  OAI31X1 g175363(.A0 (n_4819), .A1 (n_4820), .A2 (n_4994), .B0
       (cpu_state[5]), .Y (n_5087));
  AOI211XL g175364(.A0 (reg_pc[18]), .A1 (n_961), .B0 (n_4825), .C0
       (n_5016), .Y (n_5086));
  OAI2BB1X1 g175365(.A0N (n_11739), .A1N (n_5020), .B0 (n_869), .Y
       (n_5085));
  MX2X1 g175366(.A (instr_ecall_ebreak), .B (n_5014), .S0 (n_538), .Y
       (n_5084));
  AOI221X1 g175367(.A0 (\cpuregs[5] [21]), .A1 (n_11748), .B0 (n_833),
       .B1 (n_6939), .C0 (n_5038), .Y (n_5083));
  OAI32X1 g175368(.A0 (mem_rdata_q[23]), .A1 (n_537), .A2 (n_4985), .B0
       (n_709), .B1 (n_538), .Y (n_5082));
  NAND2X1 g175372(.A (n_2433), .B (n_5059), .Y (n_5098));
  AOI22X1 g175374(.A0 (mem_rdata_q[13]), .A1 (n_5025), .B0 (n_437), .B1
       (n_696), .Y (n_5081));
  AOI211XL g175375(.A0 (\cpuregs[5] [11]), .A1 (n_291), .B0 (n_4840),
       .C0 (n_5005), .Y (n_5080));
  AOI211XL g175376(.A0 (\cpuregs[5] [12]), .A1 (n_291), .B0 (n_4838),
       .C0 (n_5004), .Y (n_5079));
  AOI221X1 g175377(.A0 (\cpuregs[1] [13]), .A1 (n_456), .B0
       (\cpuregs[2] [13]), .B1 (n_425), .C0 (n_5051), .Y (n_5078));
  AOI22X1 g175378(.A0 (cpu_state[5]), .A1 (n_4995), .B0 (reg_pc[16]),
       .B1 (n_547), .Y (n_5077));
  AOI211XL g175379(.A0 (\cpuregs[5] [17]), .A1 (n_291), .B0 (n_4827),
       .C0 (n_5002), .Y (n_5076));
  AOI211XL g175380(.A0 (\cpuregs[5] [24]), .A1 (n_291), .B0 (n_4813),
       .C0 (n_5001), .Y (n_5075));
  AOI22X1 g175381(.A0 (cpu_state[5]), .A1 (n_5021), .B0 (reg_pc[25]),
       .B1 (n_547), .Y (n_5074));
  AOI221X1 g175382(.A0 (\cpuregs[1] [26]), .A1 (n_456), .B0
       (\cpuregs[2] [26]), .B1 (n_425), .C0 (n_5031), .Y (n_5073));
  AOI221X1 g175383(.A0 (\cpuregs[1] [27]), .A1 (n_456), .B0
       (\cpuregs[2] [27]), .B1 (n_425), .C0 (n_5045), .Y (n_5072));
  AOI221X1 g175384(.A0 (\cpuregs[1] [28]), .A1 (n_456), .B0
       (\cpuregs[2] [28]), .B1 (n_425), .C0 (n_5044), .Y (n_5071));
  AOI221X1 g175385(.A0 (\cpuregs[1] [29]), .A1 (n_456), .B0
       (\cpuregs[2] [29]), .B1 (n_425), .C0 (n_5043), .Y (n_5070));
  AO22X1 g175386(.A0 (n_2508), .A1 (n_5028), .B0 (cpu_state[3]), .B1
       (n_348), .Y (n_5069));
  AOI211XL g175387(.A0 (\cpuregs[15] [23]), .A1 (n_462), .B0 (n_4944),
       .C0 (n_4993), .Y (n_5068));
  OAI22X1 g175388(.A0 (n_2415), .A1 (n_5027), .B0 (n_611), .B1 (n_702),
       .Y (n_5067));
  OAI22X1 g175389(.A0 (n_973), .A1 (n_5027), .B0 (n_564), .B1 (n_702),
       .Y (n_5066));
  AOI22X1 g175390(.A0 (mem_rdata_q[28]), .A1 (n_5025), .B0 (n_2144),
       .B1 (n_14), .Y (n_5065));
  OAI22X1 g175391(.A0 (n_2334), .A1 (n_5027), .B0 (n_761), .B1 (n_702),
       .Y (n_5064));
  AOI221X1 g175392(.A0 (n_1810), .A1 (n_432), .B0 (mem_rdata_q[22]),
       .B1 (n_703), .C0 (n_3258), .Y (n_5063));
  AOI221X1 g175393(.A0 (n_2137), .A1 (n_3418), .B0 (n_440), .B1
       (n_2421), .C0 (n_5033), .Y (n_5062));
  AOI221X1 g175394(.A0 (\cpuregs[1] [10]), .A1 (n_456), .B0
       (\cpuregs[2] [10]), .B1 (n_425), .C0 (n_5050), .Y (n_5061));
  NAND4BX1 g175396(.AN (n_4845), .B (n_4504), .C (n_4505), .D (n_4984),
       .Y (n_5057));
  NAND4XL g175397(.A (n_4555), .B (n_4554), .C (n_4914), .D (n_4982),
       .Y (n_5056));
  NAND4XL g175398(.A (n_4591), .B (n_4590), .C (n_4915), .D (n_4980),
       .Y (n_5055));
  NAND2X1 g175399(.A (n_2443), .B (n_4992), .Y (n_5054));
  NAND2X1 g175400(.A (mem_rdata_q[14]), .B (n_5025), .Y (n_5053));
  NAND2X1 g175401(.A (mem_rdata_q[31]), .B (n_5025), .Y (n_5052));
  NAND3BXL g175402(.AN (n_5003), .B (n_4352), .C (n_4793), .Y (n_5051));
  NAND3BXL g175403(.AN (n_5006), .B (n_4391), .C (n_4792), .Y (n_5050));
  NAND3BXL g175404(.AN (n_5009), .B (n_4453), .C (n_4791), .Y (n_5049));
  AOI32X1 g175405(.A0 (n_4679), .A1 (n_4680), .A2 (n_4987), .B0
       (n_548), .B1 (n_1530), .Y (n_5048));
  NAND3BXL g175406(.AN (n_5011), .B (n_4520), .C (n_4789), .Y (n_5047));
  NAND2X1 g175407(.A (n_1330), .B (n_5026), .Y (n_5060));
  NOR2X1 g175408(.A (n_1590), .B (n_5025), .Y (n_5059));
  NAND2X1 g175409(.A (n_4991), .B (n_5026), .Y (n_301));
  OAI221X1 g175411(.A0 (n_682), .A1 (n_2443), .B0 (n_2145), .B1
       (n_4951), .C0 (n_1232), .Y (n_5046));
  NAND3BXL g175412(.AN (n_4999), .B (n_4649), .C (n_4753), .Y (n_5045));
  NAND3BXL g175413(.AN (n_4998), .B (n_4660), .C (n_4752), .Y (n_5044));
  NAND3BXL g175414(.AN (n_4997), .B (n_4671), .C (n_4751), .Y (n_5043));
  NAND4XL g175415(.A (mem_rdata_q[27]), .B (n_639), .C (n_977), .D
       (n_4952), .Y (n_5042));
  AOI22X1 g175416(.A0 (n_1549), .A1 (n_4989), .B0 (cpu_state[6]), .B1
       (n_348), .Y (n_5041));
  AOI221X1 g175417(.A0 (\cpuregs[1] [6]), .A1 (n_456), .B0
       (\cpuregs[2] [6]), .B1 (n_425), .C0 (n_5022), .Y (n_5040));
  AOI221X1 g175418(.A0 (\cpuregs[1] [15]), .A1 (n_456), .B0
       (\cpuregs[2] [15]), .B1 (n_425), .C0 (n_5024), .Y (n_5039));
  OAI211X1 g175419(.A0 (n_655), .A1 (n_4287), .B0 (n_4745), .C0
       (n_4981), .Y (n_5038));
  OAI22X1 g175420(.A0 (n_615), .A1 (n_4990), .B0 (n_548), .B1 (n_702),
       .Y (n_5037));
  AOI22X1 g175421(.A0 (n_1812), .A1 (n_432), .B0 (n_437), .B1 (n_2998),
       .Y (n_5036));
  AOI22X1 g175422(.A0 (n_1811), .A1 (n_432), .B0 (n_504), .B1 (n_2998),
       .Y (n_5035));
  AOI221X1 g175423(.A0 (n_687), .A1 (n_2426), .B0 (decoded_rd[0]), .B1
       (n_953), .C0 (n_4996), .Y (n_5034));
  OAI22X1 g175424(.A0 (n_1807), .A1 (n_704), .B0 (n_590), .B1 (n_341),
       .Y (n_5033));
  OAI221X1 g175425(.A0 (n_679), .A1 (n_2443), .B0 (n_2143), .B1
       (n_4951), .C0 (n_1258), .Y (n_5032));
  NAND3BXL g175426(.AN (n_5000), .B (n_4638), .C (n_4754), .Y (n_5031));
  INVX1 g175427(.A (n_5029), .Y (n_5030));
  INVX1 g175428(.A (n_5028), .Y (n_5027));
  INVX1 g175429(.A (n_5026), .Y (n_5025));
  NAND4BX1 g175430(.AN (n_4832), .B (n_4321), .C (n_4322), .D (n_4913),
       .Y (n_5024));
  NAND2X1 g175431(.A (n_1813), .B (n_432), .Y (n_5023));
  NAND4BX1 g175432(.AN (n_4870), .B (n_4437), .C (n_4438), .D (n_4911),
       .Y (n_5022));
  NOR2X1 g175433(.A (n_11691), .B (n_4962), .Y (n_5029));
  NOR2X1 g175440(.A (n_548), .B (n_4990), .Y (n_5028));
  NAND2X1 g175457(.A (n_445), .B (n_4991), .Y (n_5026));
  NAND4XL g175459(.A (n_4621), .B (n_4622), .C (n_4908), .D (n_4925),
       .Y (n_5021));
  OAI211X1 g175460(.A0 (n_6), .A1 (n_4920), .B0 (n_2113), .C0 (n_2190),
       .Y (n_5020));
  NAND4XL g175461(.A (n_1459), .B (n_4497), .C (n_4786), .D (n_4946),
       .Y (n_5019));
  NAND4XL g175462(.A (n_4483), .B (n_4484), .C (n_4785), .D (n_4947),
       .Y (n_5018));
  NAND4XL g175463(.A (n_4694), .B (n_4767), .C (n_4948), .D (n_1448),
       .Y (n_5017));
  NAND3X1 g175464(.A (n_4542), .B (n_4977), .C (n_4541), .Y (n_5016));
  NAND4XL g175465(.A (n_4342), .B (n_4779), .C (n_4949), .D (n_4343),
       .Y (n_5015));
  NOR4BX1 g175466(.AN (n_4905), .B (mem_rdata_q[7]), .C
       (mem_rdata_q[11]), .D (mem_rdata_q[10]), .Y (n_5014));
  NOR4X1 g175467(.A (\reg_op2[25]_9694 ), .B (\reg_op2[26]_9695 ), .C
       (\reg_op2[30]_9699 ), .D (n_4897), .Y (n_5013));
  OAI2BB1X1 g175468(.A0N (instr_rdcycleh), .A1N (n_537), .B0 (n_4975),
       .Y (n_5012));
  NAND4XL g175469(.A (n_4519), .B (n_4518), .C (n_4517), .D (n_4929),
       .Y (n_5011));
  NAND4XL g175470(.A (n_4462), .B (n_4463), .C (n_4461), .D (n_4937),
       .Y (n_5010));
  NAND4XL g175471(.A (n_4452), .B (n_4451), .C (n_4450), .D (n_4936),
       .Y (n_5009));
  NAND4XL g175472(.A (n_4415), .B (n_4414), .C (n_4413), .D (n_4935),
       .Y (n_5008));
  NAND4XL g175473(.A (n_4401), .B (n_4400), .C (n_4399), .D (n_4934),
       .Y (n_5007));
  NAND4XL g175474(.A (n_4390), .B (n_4389), .C (n_4388), .D (n_4933),
       .Y (n_5006));
  NAND4XL g175475(.A (n_4376), .B (n_4375), .C (n_4374), .D (n_4932),
       .Y (n_5005));
  NAND4XL g175476(.A (n_4362), .B (n_4361), .C (n_4360), .D (n_4931),
       .Y (n_5004));
  NAND4XL g175477(.A (n_4351), .B (n_4350), .C (n_4349), .D (n_4930),
       .Y (n_5003));
  NAND4XL g175478(.A (n_4294), .B (n_4295), .C (n_4293), .D (n_4928),
       .Y (n_5002));
  NAND4XL g175479(.A (n_4616), .B (n_4614), .C (n_4615), .D (n_4926),
       .Y (n_5001));
  NAND4XL g175480(.A (n_4640), .B (n_4639), .C (n_4641), .D (n_4924),
       .Y (n_5000));
  NAND4XL g175481(.A (n_4651), .B (n_4650), .C (n_4652), .D (n_4923),
       .Y (n_4999));
  NAND4XL g175482(.A (n_4661), .B (n_4662), .C (n_4663), .D (n_4922),
       .Y (n_4998));
  NAND4XL g175483(.A (n_4672), .B (n_4674), .C (n_4673), .D (n_4921),
       .Y (n_4997));
  OAI22X1 g175484(.A0 (n_689), .A1 (n_4951), .B0 (n_680), .B1 (n_2443),
       .Y (n_4996));
  NAND4XL g175485(.A (n_4315), .B (n_4316), .C (n_4909), .D (n_4938),
       .Y (n_4995));
  NAND4XL g175486(.A (n_4561), .B (n_4110), .C (n_4562), .D (n_4927),
       .Y (n_4994));
  NAND4XL g175487(.A (n_4601), .B (n_4602), .C (n_4603), .D (n_4939),
       .Y (n_4993));
  AOI221X1 g175488(.A0 (n_503), .A1 (n_316), .B0 (decoded_rd[3]), .B1
       (n_953), .C0 (n_3043), .Y (n_4992));
  INVX1 g175489(.A (n_4990), .Y (n_4989));
  NOR4X1 g175491(.A (n_4803), .B (n_4804), .C (n_4918), .D (n_4769), .Y
       (n_4987));
  OR4X1 g175492(.A (\genblk2.pcpi_div_quotient_msk [5]), .B
       (\genblk2.pcpi_div_quotient_msk [6]), .C
       (\genblk2.pcpi_div_quotient_msk [30]), .D (n_4859), .Y (n_4986));
  NAND2X1 g175493(.A (n_1343), .B (n_4952), .Y (n_4985));
  AOI221X1 g175494(.A0 (\cpuregs[4] [1]), .A1 (n_424), .B0
       (\cpuregs[5] [1]), .B1 (n_291), .C0 (n_4943), .Y (n_4984));
  AOI221X1 g175495(.A0 (\cpuregs[18] [7]), .A1 (n_492), .B0
       (\cpuregs[19] [7]), .B1 (n_502), .C0 (n_4942), .Y (n_4983));
  AOI221X1 g175496(.A0 (\cpuregs[20] [19]), .A1 (n_488), .B0
       (\cpuregs[21] [19]), .B1 (n_468), .C0 (n_4950), .Y (n_4982));
  OAI31X1 g175497(.A0 (n_4817), .A1 (n_4818), .A2 (n_4898), .B0
       (cpu_state[5]), .Y (n_4981));
  AOI221X1 g175498(.A0 (\cpuregs[8] [22]), .A1 (n_466), .B0
       (\cpuregs[7] [22]), .B1 (n_474), .C0 (n_4940), .Y (n_4980));
  OAI32X1 g175499(.A0 (n_537), .A1 (n_1342), .A2 (n_4878), .B0 (n_707),
       .B1 (n_538), .Y (n_4979));
  NAND4XL g175500(.A (n_2654), .B (n_2655), .C (n_2653), .D (n_4900),
       .Y (n_4978));
  AOI211XL g175501(.A0 (\cpuregs[4] [18]), .A1 (n_424), .B0 (n_4879),
       .C0 (n_4824), .Y (n_4977));
  AO22X1 g175502(.A0 (n_440), .A1 (n_316), .B0 (decoded_rd[4]), .B1
       (n_953), .Y (n_4976));
  NAND4XL g175503(.A (mem_rdata_q[27]), .B (n_977), .C (n_538), .D
       (n_4877), .Y (n_4975));
  NAND4XL g175504(.A (n_2167), .B (n_3044), .C (n_2533), .D (n_4799),
       .Y (n_4974));
  NAND4XL g175505(.A (n_2866), .B (n_2867), .C (n_2958), .D (n_4889),
       .Y (n_4973));
  NAND4XL g175506(.A (n_2719), .B (n_2718), .C (n_2717), .D (n_4901),
       .Y (n_4972));
  NOR2X1 g175507(.A (n_2603), .B (n_4941), .Y (n_4991));
  OR2X1 g175508(.A (n_544), .B (n_4945), .Y (n_4990));
  NOR4X1 g175509(.A (n_2421), .B (n_696), .C (n_4858), .D (n_703), .Y
       (n_432));
  NAND4XL g175510(.A (n_2780), .B (n_2781), .C (n_3049), .D (n_4887),
       .Y (n_4971));
  NAND4XL g175511(.A (n_2855), .B (n_2887), .C (n_3036), .D (n_4896),
       .Y (n_4970));
  NAND4XL g175512(.A (n_2897), .B (n_2847), .C (n_3037), .D (n_4895),
       .Y (n_4969));
  NAND4XL g175513(.A (n_2903), .B (n_2904), .C (n_3032), .D (n_4894),
       .Y (n_4968));
  NAND4XL g175514(.A (n_2946), .B (n_2945), .C (n_3031), .D (n_4893),
       .Y (n_4967));
  NAND4XL g175515(.A (n_2917), .B (n_2962), .C (n_3030), .D (n_4892),
       .Y (n_4966));
  NAND4XL g175516(.A (n_2981), .B (n_2980), .C (n_3038), .D (n_4891),
       .Y (n_4965));
  NAND4XL g175517(.A (n_2926), .B (n_2989), .C (n_3029), .D (n_4890),
       .Y (n_4964));
  NAND4XL g175518(.A (n_2815), .B (n_2816), .C (n_3059), .D (n_4902),
       .Y (n_4963));
  NAND4XL g175519(.A (n_1349), .B (n_11736), .C (n_11737), .D
       (n_11738), .Y (n_4962));
  NAND4XL g175520(.A (n_2768), .B (n_2769), .C (n_3027), .D (n_4886),
       .Y (n_4961));
  NAND4XL g175521(.A (n_2794), .B (n_2795), .C (n_3028), .D (n_4888),
       .Y (n_4960));
  NAND4XL g175522(.A (n_2755), .B (n_2756), .C (n_3050), .D (n_4885),
       .Y (n_4959));
  NAND4XL g175523(.A (n_2743), .B (n_2744), .C (n_3053), .D (n_4884),
       .Y (n_4958));
  NAND4XL g175524(.A (n_2708), .B (n_2707), .C (n_3026), .D (n_4883),
       .Y (n_4957));
  NAND4XL g175525(.A (n_2680), .B (n_2681), .C (n_3024), .D (n_4882),
       .Y (n_4956));
  NAND4XL g175526(.A (n_2643), .B (n_2644), .C (n_3057), .D (n_4881),
       .Y (n_4955));
  NAND4XL g175527(.A (n_2628), .B (n_2629), .C (n_3022), .D (n_4880),
       .Y (n_4954));
  AOI32X1 g175528(.A0 (n_503), .A1 (n_2440), .A2 (n_1620), .B0
       (mem_rdata_q[23]), .B1 (n_703), .Y (n_4953));
  NAND3BXL g175529(.AN (n_4822), .B (n_4111), .C (n_4556), .Y (n_4950));
  NOR4X1 g175530(.A (n_4112), .B (n_4835), .C (n_4833), .D (n_4834), .Y
       (n_4949));
  NOR4X1 g175531(.A (n_4106), .B (n_4802), .C (n_4801), .D (n_4800), .Y
       (n_4948));
  NOR4X1 g175532(.A (n_4115), .B (n_4864), .C (n_4865), .D (n_4866), .Y
       (n_4947));
  NOR4X1 g175533(.A (n_4116), .B (n_4863), .C (n_4862), .D (n_4861), .Y
       (n_4946));
  AOI22X1 g175534(.A0 (n_975), .A1 (n_702), .B0 (n_1351), .B1 (n_4288),
       .Y (n_4945));
  OAI2BB1X1 g175535(.A0N (\cpuregs[1] [23]), .A1N (n_456), .B0
       (n_4916), .Y (n_4944));
  NAND3BXL g175536(.AN (n_4860), .B (n_4117), .C (n_4503), .Y (n_4943));
  NAND3BXL g175537(.AN (n_4873), .B (n_4113), .C (n_4427), .Y (n_4942));
  OAI221X1 g175538(.A0 (n_1329), .A1 (n_4766), .B0 (n_3005), .B1
       (n_1590), .C0 (n_3007), .Y (n_4941));
  NAND3BXL g175539(.AN (n_4815), .B (n_4109), .C (n_4592), .Y (n_4940));
  AOI221X1 g175540(.A0 (\cpuregs[22] [23]), .A1 (n_482), .B0
       (\cpuregs[23] [23]), .B1 (n_464), .C0 (n_4917), .Y (n_4939));
  NOR4X1 g175542(.A (mem_rdata_q[22]), .B (mem_rdata_q[20]), .C
       (n_644), .D (n_306), .Y (n_4952));
  NOR2X1 g175544(.A (n_3043), .B (n_316), .Y (n_4951));
  AOI221X1 g175548(.A0 (\cpuregs[1] [16]), .A1 (n_456), .B0
       (\cpuregs[3] [16]), .B1 (n_423), .C0 (n_4830), .Y (n_4938));
  AOI221X1 g175549(.A0 (\cpuregs[26] [4]), .A1 (n_490), .B0
       (\cpuregs[29] [4]), .B1 (n_458), .C0 (n_4868), .Y (n_4937));
  AOI221X1 g175550(.A0 (\cpuregs[18] [5]), .A1 (n_492), .B0
       (\cpuregs[21] [5]), .B1 (n_468), .C0 (n_4869), .Y (n_4936));
  AOI221X1 g175551(.A0 (\cpuregs[22] [8]), .A1 (n_482), .B0
       (\cpuregs[19] [8]), .B1 (n_502), .C0 (n_4875), .Y (n_4935));
  AOI221X1 g175552(.A0 (\cpuregs[22] [9]), .A1 (n_482), .B0
       (\cpuregs[21] [9]), .B1 (n_468), .C0 (n_4842), .Y (n_4934));
  AOI221X1 g175553(.A0 (\cpuregs[24] [10]), .A1 (n_494), .B0
       (\cpuregs[31] [10]), .B1 (n_476), .C0 (n_4841), .Y (n_4933));
  AOI221X1 g175554(.A0 (\cpuregs[18] [11]), .A1 (n_492), .B0
       (\cpuregs[23] [11]), .B1 (n_464), .C0 (n_4839), .Y (n_4932));
  AOI221X1 g175555(.A0 (\cpuregs[26] [12]), .A1 (n_490), .B0
       (\cpuregs[29] [12]), .B1 (n_458), .C0 (n_4837), .Y (n_4931));
  AOI221X1 g175556(.A0 (\cpuregs[24] [13]), .A1 (n_494), .B0
       (\cpuregs[31] [13]), .B1 (n_476), .C0 (n_4836), .Y (n_4930));
  AOI221X1 g175557(.A0 (\cpuregs[22] [0]), .A1 (n_482), .B0
       (\cpuregs[17] [0]), .B1 (n_486), .C0 (n_4844), .Y (n_4929));
  AOI221X1 g175558(.A0 (\cpuregs[26] [17]), .A1 (n_490), .B0
       (\cpuregs[31] [17]), .B1 (n_476), .C0 (n_4826), .Y (n_4928));
  AOI221X1 g175559(.A0 (\cpuregs[15] [20]), .A1 (n_462), .B0
       (\cpuregs[5] [20]), .B1 (n_291), .C0 (n_4821), .Y (n_4927));
  AOI221X1 g175560(.A0 (\cpuregs[26] [24]), .A1 (n_490), .B0
       (\cpuregs[31] [24]), .B1 (n_476), .C0 (n_4812), .Y (n_4926));
  AOI221X1 g175561(.A0 (\cpuregs[5] [25]), .A1 (n_291), .B0
       (\cpuregs[15] [25]), .B1 (n_462), .C0 (n_4811), .Y (n_4925));
  AOI221X1 g175562(.A0 (\cpuregs[26] [26]), .A1 (n_490), .B0
       (\cpuregs[29] [26]), .B1 (n_458), .C0 (n_4808), .Y (n_4924));
  AOI221X1 g175563(.A0 (\cpuregs[26] [27]), .A1 (n_490), .B0
       (\cpuregs[29] [27]), .B1 (n_458), .C0 (n_4807), .Y (n_4923));
  AOI221X1 g175564(.A0 (\cpuregs[22] [28]), .A1 (n_482), .B0
       (\cpuregs[21] [28]), .B1 (n_468), .C0 (n_4806), .Y (n_4922));
  AOI221X1 g175565(.A0 (\cpuregs[24] [29]), .A1 (n_494), .B0
       (\cpuregs[27] [29]), .B1 (n_498), .C0 (n_4805), .Y (n_4921));
  OAI211X1 g175566(.A0 (n_856), .A1 (n_4775), .B0 (n_884), .C0 (n_863),
       .Y (n_4920));
  OAI211X1 g175567(.A0 (n_611), .A1 (n_1903), .B0 (n_2165), .C0
       (n_4737), .Y (n_4919));
  NAND4XL g175568(.A (n_4107), .B (n_4684), .C (n_4683), .D (n_4768),
       .Y (n_4918));
  NAND4XL g175569(.A (n_4108), .B (n_4606), .C (n_4605), .D (n_4774),
       .Y (n_4917));
  AOI221X1 g175570(.A0 (\cpuregs[4] [23]), .A1 (n_424), .B0
       (\cpuregs[3] [23]), .B1 (n_423), .C0 (n_4814), .Y (n_4916));
  AOI221X1 g175571(.A0 (\cpuregs[1] [22]), .A1 (n_456), .B0
       (\cpuregs[15] [22]), .B1 (n_462), .C0 (n_4816), .Y (n_4915));
  AOI221X1 g175572(.A0 (\cpuregs[2] [19]), .A1 (n_425), .B0
       (\cpuregs[15] [19]), .B1 (n_462), .C0 (n_4823), .Y (n_4914));
  AOI21X1 g175573(.A0 (\cpuregs[15] [15]), .A1 (n_462), .B0 (n_4831),
       .Y (n_4913));
  AOI221X1 g175574(.A0 (\cpuregs[4] [7]), .A1 (n_424), .B0
       (\cpuregs[3] [7]), .B1 (n_423), .C0 (n_4872), .Y (n_4912));
  AOI21X1 g175575(.A0 (\cpuregs[15] [6]), .A1 (n_462), .B0 (n_4871), .Y
       (n_4911));
  NAND3BXL g175576(.AN (n_3043), .B (n_2511), .C (n_4757), .Y (n_4910));
  NOR2X1 g175577(.A (n_4828), .B (n_4829), .Y (n_4909));
  NOR2X1 g175578(.A (n_4809), .B (n_4810), .Y (n_4908));
  OAI211X1 g175579(.A0 (n_2143), .A1 (n_296), .B0 (n_1299), .C0
       (n_2168), .Y (n_4907));
  OAI211X1 g175580(.A0 (n_611), .A1 (n_16), .B0 (n_2165), .C0 (n_4736),
       .Y (n_4906));
  AOI211XL g175581(.A0 (n_2479), .A1 (n_4529), .B0 (mem_rdata_q[8]),
       .C0 (mem_rdata_q[9]), .Y (n_4905));
  AOI211XL g175593(.A0 (\cpuregs[14] [16]), .A1 (n_2531), .B0 (n_3134),
       .C0 (n_4725), .Y (n_4902));
  AOI221X1 g175594(.A0 (\cpuregs[24] [24]), .A1 (n_2490), .B0
       (\cpuregs[23] [24]), .B1 (n_2500), .C0 (n_4797), .Y (n_4901));
  AOI221X1 g175595(.A0 (\cpuregs[28] [29]), .A1 (n_2491), .B0
       (\cpuregs[27] [29]), .B1 (n_2525), .C0 (n_4796), .Y (n_4900));
  OAI211X1 g175596(.A0 (n_689), .A1 (n_296), .B0 (n_1282), .C0
       (n_2335), .Y (n_4899));
  NAND4XL g175597(.A (n_4575), .B (n_4576), .C (n_4776), .D (n_4755),
       .Y (n_4898));
  NAND4XL g175598(.A (\genblk2.pcpi_div_minus_2470_59_n_474 ), .B
       (n_746), .C (n_630), .D (n_4530), .Y (n_4897));
  AOI211XL g175599(.A0 (\cpuregs[14] [8]), .A1 (n_2531), .B0 (n_3123),
       .C0 (n_4732), .Y (n_4896));
  AOI211XL g175600(.A0 (\cpuregs[14] [9]), .A1 (n_2531), .B0 (n_3122),
       .C0 (n_4731), .Y (n_4895));
  AOI211XL g175601(.A0 (\cpuregs[14] [11]), .A1 (n_2531), .B0 (n_3117),
       .C0 (n_4730), .Y (n_4894));
  AOI211XL g175602(.A0 (\cpuregs[14] [12]), .A1 (n_2531), .B0 (n_3132),
       .C0 (n_4729), .Y (n_4893));
  AOI211XL g175603(.A0 (\cpuregs[14] [13]), .A1 (n_2531), .B0 (n_3115),
       .C0 (n_4728), .Y (n_4892));
  AOI211XL g175604(.A0 (\cpuregs[14] [14]), .A1 (n_2531), .B0 (n_3113),
       .C0 (n_4727), .Y (n_4891));
  AOI211XL g175605(.A0 (\cpuregs[14] [15]), .A1 (n_2531), .B0 (n_3111),
       .C0 (n_4726), .Y (n_4890));
  AOI221X1 g175606(.A0 (\cpuregs[29] [7]), .A1 (n_2524), .B0
       (\cpuregs[30] [7]), .B1 (n_2523), .C0 (n_4798), .Y (n_4889));
  AOI211XL g175607(.A0 (\cpuregs[14] [18]), .A1 (n_2531), .B0 (n_3104),
       .C0 (n_4724), .Y (n_4888));
  AOI211XL g175608(.A0 (\cpuregs[14] [19]), .A1 (n_2531), .B0 (n_3102),
       .C0 (n_4723), .Y (n_4887));
  AOI211XL g175609(.A0 (\cpuregs[14] [20]), .A1 (n_2531), .B0 (n_3100),
       .C0 (n_4722), .Y (n_4886));
  AOI211XL g175610(.A0 (\cpuregs[14] [21]), .A1 (n_2531), .B0 (n_3098),
       .C0 (n_4721), .Y (n_4885));
  AOI211XL g175611(.A0 (\cpuregs[14] [22]), .A1 (n_2531), .B0 (n_3096),
       .C0 (n_4720), .Y (n_4884));
  AOI211XL g175612(.A0 (\cpuregs[14] [25]), .A1 (n_2531), .B0 (n_3090),
       .C0 (n_4719), .Y (n_4883));
  AOI211XL g175613(.A0 (\cpuregs[14] [27]), .A1 (n_2531), .B0 (n_3085),
       .C0 (n_4718), .Y (n_4882));
  AOI211XL g175614(.A0 (\cpuregs[14] [30]), .A1 (n_2531), .B0 (n_3080),
       .C0 (n_4717), .Y (n_4881));
  AOI211XL g175615(.A0 (\cpuregs[14] [31]), .A1 (n_2531), .B0 (n_3078),
       .C0 (n_4716), .Y (n_4880));
  NAND4XL g175616(.A (n_4549), .B (n_4548), .C (n_4713), .D (n_4777),
       .Y (n_4879));
  NAND3BXL g175617(.AN (n_4756), .B (n_342), .C (n_3044), .Y (n_316));
  NAND4XL g175618(.A (n_445), .B (n_2606), .C (n_4712), .D (n_3007), .Y
       (n_341));
  INVX1 g175619(.A (n_4877), .Y (n_4878));
  NAND4XL g175621(.A (n_4409), .B (n_4412), .C (n_4411), .D (n_4410),
       .Y (n_4875));
  NAND4XL g175622(.A (n_4419), .B (n_4418), .C (n_4417), .D (n_4416),
       .Y (n_4874));
  NAND4XL g175623(.A (n_4423), .B (n_4426), .C (n_4425), .D (n_4424),
       .Y (n_4873));
  NAND4XL g175624(.A (n_4429), .B (n_4431), .C (n_4432), .D (n_4430),
       .Y (n_4872));
  NAND4XL g175625(.A (n_4433), .B (n_4435), .C (n_4436), .D (n_4434),
       .Y (n_4871));
  NAND4XL g175626(.A (n_4439), .B (n_4442), .C (n_4441), .D (n_4440),
       .Y (n_4870));
  NAND4XL g175627(.A (n_4446), .B (n_4449), .C (n_4448), .D (n_4447),
       .Y (n_4869));
  NAND4XL g175628(.A (n_4457), .B (n_4460), .C (n_4459), .D (n_4458),
       .Y (n_4868));
  NAND4XL g175629(.A (n_4467), .B (n_4464), .C (n_4466), .D (n_4465),
       .Y (n_4867));
  NAND4XL g175630(.A (n_4475), .B (n_4478), .C (n_4477), .D (n_4476),
       .Y (n_4866));
  NAND4XL g175631(.A (n_4471), .B (n_4474), .C (n_4473), .D (n_4472),
       .Y (n_4865));
  NAND4XL g175632(.A (n_4482), .B (n_4479), .C (n_4481), .D (n_4480),
       .Y (n_4864));
  NAND4XL g175633(.A (n_4485), .B (n_4488), .C (n_4487), .D (n_4486),
       .Y (n_4863));
  NAND4XL g175634(.A (n_4489), .B (n_4492), .C (n_4491), .D (n_4490),
       .Y (n_4862));
  NAND4XL g175635(.A (n_4493), .B (n_4496), .C (n_4495), .D (n_4494),
       .Y (n_4861));
  NAND4XL g175636(.A (n_4500), .B (n_4499), .C (n_4502), .D (n_4501),
       .Y (n_4860));
  OR4X1 g175637(.A (\genblk2.pcpi_div_quotient_msk [29]), .B
       (\genblk2.pcpi_div_quotient_msk [28]), .C
       (\genblk2.pcpi_div_quotient_msk [27]), .D (n_4105), .Y (n_4859));
  NAND3BXL g175638(.AN (n_2998), .B (n_4712), .C (n_3065), .Y (n_4858));
  AOI221X1 g175639(.A0 (\cpuregs[5] [19]), .A1 (n_11748), .B0 (n_833),
       .B1 (n_6941), .C0 (n_4747), .Y (n_4857));
  AOI221X1 g175640(.A0 (\cpuregs[5] [22]), .A1 (n_11748), .B0 (n_833),
       .B1 (n_6938), .C0 (n_4744), .Y (n_4856));
  OAI211X1 g175641(.A0 (n_643), .A1 (n_35), .B0 (n_2535), .C0 (n_4533),
       .Y (n_4855));
  OAI211X1 g175642(.A0 (n_633), .A1 (n_969), .B0 (n_2111), .C0
       (n_4535), .Y (n_4854));
  OAI222X1 g175643(.A0 (n_647), .A1 (n_35), .B0 (n_2145), .B1 (n_4290),
       .C0 (n_682), .C1 (n_2437), .Y (n_4853));
  OAI2BB1X1 g175644(.A0N (decoded_imm[0]), .A1N (n_421), .B0 (n_4740),
       .Y (n_4852));
  OAI2BB1X1 g175645(.A0N (decoded_imm[1]), .A1N (n_421), .B0 (n_4739),
       .Y (n_4851));
  OAI2BB1X1 g175646(.A0N (decoded_imm[4]), .A1N (n_421), .B0 (n_4738),
       .Y (n_4850));
  OAI211X1 g175647(.A0 (n_682), .A1 (n_349), .B0 (n_1304), .C0
       (n_2171), .Y (n_4849));
  OAI211X1 g175648(.A0 (n_679), .A1 (n_349), .B0 (n_1303), .C0
       (n_2172), .Y (n_4848));
  OAI221X1 g175649(.A0 (n_680), .A1 (n_349), .B0 (n_633), .B1 (n_667),
       .C0 (n_2173), .Y (n_4847));
  NAND4XL g175650(.A (n_3250), .B (n_2584), .C (n_2605), .D (n_3495),
       .Y (n_4846));
  NAND4XL g175651(.A (n_4506), .B (n_4509), .C (n_4508), .D (n_4507),
       .Y (n_4845));
  NAND4XL g175652(.A (n_4513), .B (n_4516), .C (n_4515), .D (n_4514),
       .Y (n_4844));
  NOR2BX1 g175653(.AN (n_1356), .B (n_306), .Y (n_4877));
  NOR4X1 g175666(.A (n_849), .B (n_544), .C (n_303), .D (n_4288), .Y
       (n_348));
  NAND4XL g175671(.A (n_4395), .B (n_4398), .C (n_4397), .D (n_4396),
       .Y (n_4842));
  NAND4XL g175672(.A (n_4384), .B (n_4387), .C (n_4386), .D (n_4385),
       .Y (n_4841));
  NAND4XL g175673(.A (n_4379), .B (n_4380), .C (n_4378), .D (n_4377),
       .Y (n_4840));
  NAND4XL g175674(.A (n_4370), .B (n_4373), .C (n_4372), .D (n_4371),
       .Y (n_4839));
  NAND4XL g175675(.A (n_4363), .B (n_4366), .C (n_4365), .D (n_4364),
       .Y (n_4838));
  NAND4XL g175676(.A (n_4356), .B (n_4359), .C (n_4358), .D (n_4357),
       .Y (n_4837));
  NAND4XL g175677(.A (n_4345), .B (n_4348), .C (n_4347), .D (n_4346),
       .Y (n_4836));
  NAND4XL g175678(.A (n_4341), .B (n_4338), .C (n_4340), .D (n_4339),
       .Y (n_4835));
  NAND4XL g175679(.A (n_4334), .B (n_4337), .C (n_4336), .D (n_4335),
       .Y (n_4834));
  NAND4XL g175680(.A (n_4330), .B (n_4333), .C (n_4332), .D (n_4331),
       .Y (n_4833));
  NAND4XL g175681(.A (n_4323), .B (n_4326), .C (n_4325), .D (n_4324),
       .Y (n_4832));
  NAND4XL g175682(.A (n_4320), .B (n_4317), .C (n_4319), .D (n_4318),
       .Y (n_4831));
  NAND4XL g175683(.A (n_4312), .B (n_4314), .C (n_4311), .D (n_4313),
       .Y (n_4830));
  NAND4XL g175684(.A (n_4307), .B (n_4310), .C (n_4309), .D (n_4308),
       .Y (n_4829));
  NAND4XL g175685(.A (n_4303), .B (n_4306), .C (n_4305), .D (n_4304),
       .Y (n_4828));
  NAND4XL g175686(.A (n_4299), .B (n_4298), .C (n_4297), .D (n_4296),
       .Y (n_4827));
  NAND4XL g175687(.A (n_4536), .B (n_4292), .C (n_4291), .D (n_4531),
       .Y (n_4826));
  NAND4XL g175688(.A (n_4540), .B (n_4538), .C (n_4537), .D (n_4539),
       .Y (n_4825));
  NAND4XL g175689(.A (n_4546), .B (n_4544), .C (n_4545), .D (n_4543),
       .Y (n_4824));
  NAND4XL g175690(.A (n_4550), .B (n_4553), .C (n_4551), .D (n_4552),
       .Y (n_4823));
  NAND4XL g175691(.A (n_4560), .B (n_4557), .C (n_4558), .D (n_4559),
       .Y (n_4822));
  NAND4XL g175692(.A (n_4566), .B (n_4563), .C (n_4564), .D (n_4565),
       .Y (n_4821));
  NAND4XL g175693(.A (n_4570), .B (n_4567), .C (n_4568), .D (n_4569),
       .Y (n_4820));
  NAND4XL g175694(.A (n_4574), .B (n_4571), .C (n_4572), .D (n_4573),
       .Y (n_4819));
  NAND4XL g175695(.A (n_4581), .B (n_4578), .C (n_4579), .D (n_4580),
       .Y (n_4818));
  NAND4XL g175696(.A (n_4585), .B (n_4583), .C (n_4584), .D (n_4582),
       .Y (n_4817));
  NAND4XL g175697(.A (n_4589), .B (n_4586), .C (n_4587), .D (n_4588),
       .Y (n_4816));
  NAND4XL g175698(.A (n_4595), .B (n_4593), .C (n_4594), .D (n_4596),
       .Y (n_4815));
  NAND4XL g175699(.A (n_4600), .B (n_4597), .C (n_4598), .D (n_4599),
       .Y (n_4814));
  NAND4XL g175700(.A (n_4612), .B (n_4610), .C (n_4613), .D (n_4611),
       .Y (n_4813));
  NAND4XL g175701(.A (n_4620), .B (n_4617), .C (n_4618), .D (n_4619),
       .Y (n_4812));
  NAND4XL g175702(.A (n_4625), .B (n_4623), .C (n_4626), .D (n_4624),
       .Y (n_4811));
  NAND4XL g175703(.A (n_4630), .B (n_4627), .C (n_4628), .D (n_4629),
       .Y (n_4810));
  NAND4XL g175704(.A (n_4634), .B (n_4631), .C (n_4632), .D (n_4633),
       .Y (n_4809));
  NAND4XL g175705(.A (n_4645), .B (n_4642), .C (n_4643), .D (n_4644),
       .Y (n_4808));
  NAND4XL g175706(.A (n_4656), .B (n_4653), .C (n_4654), .D (n_4655),
       .Y (n_4807));
  NAND4XL g175707(.A (n_4667), .B (n_4664), .C (n_4665), .D (n_4666),
       .Y (n_4806));
  NAND4XL g175708(.A (n_4678), .B (n_4675), .C (n_4676), .D (n_4677),
       .Y (n_4805));
  NAND4XL g175709(.A (n_4688), .B (n_4685), .C (n_4686), .D (n_4687),
       .Y (n_4804));
  NAND4XL g175710(.A (n_4692), .B (n_4689), .C (n_4690), .D (n_4691),
       .Y (n_4803));
  NAND4XL g175711(.A (n_4697), .B (n_4695), .C (n_4698), .D (n_4696),
       .Y (n_4802));
  NAND4XL g175712(.A (n_4706), .B (n_4703), .C (n_4704), .D (n_4705),
       .Y (n_4801));
  NAND4XL g175713(.A (n_4702), .B (n_4699), .C (n_4700), .D (n_4701),
       .Y (n_4800));
  AOI221X1 g175714(.A0 (n_2435), .A1 (n_1619), .B0 (decoded_rs1[1]),
       .B1 (n_953), .C0 (n_4788), .Y (n_4799));
  NAND4XL g175715(.A (n_1538), .B (n_2862), .C (n_2863), .D (n_4526),
       .Y (n_4798));
  NAND4XL g175716(.A (n_1539), .B (n_2715), .C (n_2716), .D (n_4525),
       .Y (n_4797));
  NAND4XL g175717(.A (n_1527), .B (n_2651), .C (n_2652), .D (n_4524),
       .Y (n_4796));
  NAND4XL g175718(.A (n_4404), .B (n_4405), .C (n_4403), .D (n_4402),
       .Y (n_4795));
  AOI221X1 g175719(.A0 (\cpuregs[12] [26]), .A1 (n_484), .B0
       (\cpuregs[13] [26]), .B1 (n_454), .C0 (n_4637), .Y (n_4794));
  AOI222X1 g175720(.A0 (\cpuregs[4] [13]), .A1 (n_424), .B0
       (\cpuregs[5] [13]), .B1 (n_291), .C0 (\cpuregs[15] [13]), .C1
       (n_462), .Y (n_4793));
  AOI222X1 g175721(.A0 (\cpuregs[6] [10]), .A1 (n_333), .B0
       (\cpuregs[4] [10]), .B1 (n_424), .C0 (\cpuregs[15] [10]), .C1
       (n_462), .Y (n_4792));
  AOI222X1 g175722(.A0 (\cpuregs[5] [5]), .A1 (n_291), .B0
       (\cpuregs[3] [5]), .B1 (n_423), .C0 (\cpuregs[15] [5]), .C1
       (n_462), .Y (n_4791));
  NAND2X1 g175723(.A (n_4709), .B (n_3045), .Y (n_4790));
  AOI222X1 g175724(.A0 (\cpuregs[4] [0]), .A1 (n_424), .B0
       (\cpuregs[5] [0]), .B1 (n_291), .C0 (\cpuregs[15] [0]), .C1
       (n_462), .Y (n_4789));
  NOR2X1 g175725(.A (n_2145), .B (n_296), .Y (n_4788));
  AOI221X1 g175726(.A0 (\cpuregs[12] [0]), .A1 (n_484), .B0
       (\cpuregs[13] [0]), .B1 (n_454), .C0 (n_4521), .Y (n_4787));
  AOI221X1 g175727(.A0 (\cpuregs[4] [2]), .A1 (n_424), .B0
       (\cpuregs[3] [2]), .B1 (n_423), .C0 (n_4498), .Y (n_4786));
  AOI221X1 g175728(.A0 (\cpuregs[2] [3]), .A1 (n_425), .B0
       (\cpuregs[15] [3]), .B1 (n_462), .C0 (n_1458), .Y (n_4785));
  AOI221X1 g175729(.A0 (\cpuregs[10] [5]), .A1 (n_452), .B0
       (\cpuregs[7] [5]), .B1 (n_474), .C0 (n_4454), .Y (n_4784));
  AOI221X1 g175730(.A0 (\cpuregs[22] [6]), .A1 (n_482), .B0
       (\cpuregs[23] [6]), .B1 (n_464), .C0 (n_4443), .Y (n_4783));
  AOI221X1 g175731(.A0 (\cpuregs[16] [7]), .A1 (n_478), .B0
       (\cpuregs[17] [7]), .B1 (n_486), .C0 (n_4428), .Y (n_4782));
  AOI221X1 g175732(.A0 (\cpuregs[12] [10]), .A1 (n_484), .B0
       (\cpuregs[13] [10]), .B1 (n_454), .C0 (n_4392), .Y (n_4781));
  AOI221X1 g175733(.A0 (\cpuregs[7] [13]), .A1 (n_474), .B0
       (\cpuregs[11] [13]), .B1 (n_448), .C0 (n_4353), .Y (n_4780));
  AOI221X1 g175734(.A0 (\cpuregs[3] [14]), .A1 (n_423), .B0
       (\cpuregs[6] [14]), .B1 (n_333), .C0 (n_4344), .Y (n_4779));
  AOI221X1 g175735(.A0 (\cpuregs[18] [15]), .A1 (n_492), .B0
       (\cpuregs[19] [15]), .B1 (n_502), .C0 (n_4327), .Y (n_4778));
  AOI221X1 g175736(.A0 (\cpuregs[9] [18]), .A1 (n_470), .B0
       (\cpuregs[7] [18]), .B1 (n_474), .C0 (n_4547), .Y (n_4777));
  AOI221X1 g175737(.A0 (\cpuregs[1] [21]), .A1 (n_456), .B0
       (\cpuregs[9] [21]), .B1 (n_470), .C0 (n_4577), .Y (n_4776));
  AOI31X1 g175738(.A0 (n_870), .A1 (n_6536), .A2 (n_3425), .B0 (n_873),
       .Y (n_4775));
  AOI221X1 g175739(.A0 (\cpuregs[26] [23]), .A1 (n_490), .B0
       (\cpuregs[27] [23]), .B1 (n_498), .C0 (n_4604), .Y (n_4774));
  OAI221X1 g175740(.A0 (n_1958), .A1 (n_3465), .B0 (n_728), .B1
       (n_3236), .C0 (n_329), .Y (n_4773));
  AOI221X1 g175741(.A0 (\cpuregs[12] [27]), .A1 (n_484), .B0
       (\cpuregs[13] [27]), .B1 (n_454), .C0 (n_4648), .Y (n_4772));
  AOI221X1 g175742(.A0 (\cpuregs[9] [28]), .A1 (n_470), .B0
       (\cpuregs[12] [28]), .B1 (n_484), .C0 (n_4659), .Y (n_4771));
  AOI221X1 g175743(.A0 (\cpuregs[8] [29]), .A1 (n_466), .B0
       (\cpuregs[7] [29]), .B1 (n_474), .C0 (n_4668), .Y (n_4770));
  NAND2X1 g175744(.A (n_4681), .B (n_1467), .Y (n_4769));
  AOI221X1 g175745(.A0 (\cpuregs[12] [30]), .A1 (n_484), .B0
       (\cpuregs[13] [30]), .B1 (n_454), .C0 (n_4682), .Y (n_4768));
  AOI221X1 g175746(.A0 (\cpuregs[4] [31]), .A1 (n_424), .B0
       (\cpuregs[3] [31]), .B1 (n_423), .C0 (n_4693), .Y (n_4767));
  NOR4X1 g175747(.A (n_2318), .B (n_2317), .C (n_2955), .D (n_1), .Y
       (n_4766));
  NAND4XL g175748(.A (n_2919), .B (n_2891), .C (n_3035), .D (n_4092),
       .Y (n_4765));
  NAND4XL g175749(.A (n_2877), .B (n_2878), .C (n_3034), .D (n_4091),
       .Y (n_4764));
  NAND4XL g175750(.A (n_2837), .B (n_2912), .C (n_3033), .D (n_4090),
       .Y (n_4763));
  NAND4XL g175751(.A (n_2806), .B (n_2807), .C (n_3058), .D (n_4089),
       .Y (n_4762));
  NAND4XL g175752(.A (n_2730), .B (n_2731), .C (n_3054), .D (n_4088),
       .Y (n_4761));
  NAND4XL g175753(.A (n_2694), .B (n_2695), .C (n_3025), .D (n_4087),
       .Y (n_4760));
  NAND4XL g175754(.A (n_2668), .B (n_2669), .C (n_3023), .D (n_4086),
       .Y (n_4759));
  NAND3BXL g175755(.AN (n_2175), .B (n_2602), .C (n_4083), .Y (n_4758));
  AOI221X1 g175756(.A0 (n_503), .A1 (n_3466), .B0 (decoded_rs1[3]), .B1
       (n_953), .C0 (n_2169), .Y (n_4757));
  OAI211X1 g175762(.A0 (n_327), .A1 (n_3412), .B0 (n_2584), .C0
       (n_3008), .Y (n_4756));
  AOI222X1 g175763(.A0 (\cpuregs[7] [21]), .A1 (n_474), .B0
       (\cpuregs[2] [21]), .B1 (n_425), .C0 (\cpuregs[15] [21]), .C1
       (n_462), .Y (n_4755));
  AOI222X1 g175764(.A0 (\cpuregs[6] [26]), .A1 (n_333), .B0
       (\cpuregs[3] [26]), .B1 (n_423), .C0 (\cpuregs[15] [26]), .C1
       (n_462), .Y (n_4754));
  AOI222X1 g175765(.A0 (\cpuregs[4] [27]), .A1 (n_424), .B0
       (\cpuregs[5] [27]), .B1 (n_291), .C0 (\cpuregs[15] [27]), .C1
       (n_462), .Y (n_4753));
  AOI222X1 g175766(.A0 (\cpuregs[3] [28]), .A1 (n_423), .B0
       (\cpuregs[5] [28]), .B1 (n_291), .C0 (\cpuregs[15] [28]), .C1
       (n_462), .Y (n_4752));
  AOI222X1 g175767(.A0 (\cpuregs[6] [29]), .A1 (n_333), .B0
       (\cpuregs[3] [29]), .B1 (n_423), .C0 (\cpuregs[15] [29]), .C1
       (n_462), .Y (n_4751));
  AOI22X1 g175768(.A0 (\cpuregs[6] [7]), .A1 (n_11746), .B0
       (\reg_op1[3]_9640 ), .B1 (n_1944), .Y (n_4750));
  AOI22X1 g175769(.A0 (\cpuregs[2] [7]), .A1 (n_11743), .B0
       (\cpuregs[5] [7]), .B1 (n_11748), .Y (n_4749));
  AOI22X1 g175770(.A0 (\cpuregs[2] [16]), .A1 (n_11743), .B0
       (\reg_op1[17]_9654 ), .B1 (n_550), .Y (n_4748));
  AO22X1 g175771(.A0 (\cpuregs[4] [19]), .A1 (n_11744), .B0
       (\cpuregs[6] [19]), .B1 (n_11746), .Y (n_4747));
  OAI22X1 g175772(.A0 (n_604), .A1 (n_4287), .B0 (n_619), .B1 (n_1943),
       .Y (n_4746));
  AOI22X1 g175773(.A0 (\cpuregs[4] [21]), .A1 (n_11744), .B0
       (\cpuregs[6] [21]), .B1 (n_11746), .Y (n_4745));
  AO22X1 g175774(.A0 (\cpuregs[4] [22]), .A1 (n_11744), .B0
       (\cpuregs[6] [22]), .B1 (n_11746), .Y (n_4744));
  OAI22X1 g175775(.A0 (n_606), .A1 (n_4287), .B0 (n_625), .B1 (n_1943),
       .Y (n_4743));
  AOI22X1 g175776(.A0 (\cpuregs[6] [23]), .A1 (n_11746), .B0
       (\reg_op1[19]_9656 ), .B1 (n_1944), .Y (n_4742));
  AOI22X1 g175777(.A0 (\cpuregs[2] [25]), .A1 (n_11743), .B0
       (\reg_op1[26]_9663 ), .B1 (n_550), .Y (n_4741));
  AOI22X1 g175778(.A0 (n_310), .A1 (n_344), .B0 (\reg_op2[0]_9669 ),
       .B1 (n_832), .Y (n_4740));
  AOI22X1 g175779(.A0 (n_309), .A1 (n_344), .B0 (\reg_op2[1]_9670 ),
       .B1 (n_832), .Y (n_4739));
  AOI22X1 g175780(.A0 (n_300), .A1 (n_344), .B0 (\reg_op2[4]_9673 ),
       .B1 (n_832), .Y (n_4738));
  AOI22X1 g175781(.A0 (n_2441), .A1 (n_309), .B0 (decoded_rs2[1]), .B1
       (n_968), .Y (n_4737));
  AOI22X1 g175782(.A0 (n_2441), .A1 (n_300), .B0 (decoded_rs2[4]), .B1
       (n_968), .Y (n_4736));
  OAI221X1 g175783(.A0 (n_1815), .A1 (n_3465), .B0 (n_597), .B1
       (n_3236), .C0 (n_329), .Y (n_4735));
  OAI211X1 g175784(.A0 (n_574), .A1 (n_667), .B0 (n_2176), .C0
       (n_4104), .Y (n_4734));
  OAI221X1 g175785(.A0 (n_1803), .A1 (n_3465), .B0 (n_596), .B1
       (n_3236), .C0 (n_329), .Y (n_4733));
  NAND4XL g175786(.A (n_2851), .B (n_2850), .C (n_2993), .D (n_3489),
       .Y (n_4732));
  NAND4XL g175787(.A (n_2844), .B (n_2843), .C (n_2842), .D (n_3488),
       .Y (n_4731));
  NAND4XL g175788(.A (n_2906), .B (n_2825), .C (n_2824), .D (n_3487),
       .Y (n_4730));
  NAND4XL g175789(.A (n_2956), .B (n_2957), .C (n_2914), .D (n_3486),
       .Y (n_4729));
  NAND4XL g175790(.A (n_2974), .B (n_2975), .C (n_2976), .D (n_3485),
       .Y (n_4728));
  NAND4XL g175791(.A (n_2984), .B (n_2923), .C (n_2924), .D (n_3484),
       .Y (n_4727));
  NAND4XL g175792(.A (n_2714), .B (n_2820), .C (n_2819), .D (n_3483),
       .Y (n_4726));
  NAND4XL g175793(.A (n_2810), .B (n_2936), .C (n_2937), .D (n_3482),
       .Y (n_4725));
  NAND4XL g175794(.A (n_2789), .B (n_2788), .C (n_2787), .D (n_3481),
       .Y (n_4724));
  NAND4XL g175795(.A (n_2776), .B (n_2775), .C (n_2774), .D (n_3480),
       .Y (n_4723));
  NAND4XL g175796(.A (n_2762), .B (n_2763), .C (n_2761), .D (n_3479),
       .Y (n_4722));
  NAND4XL g175797(.A (n_2751), .B (n_2750), .C (n_2749), .D (n_3478),
       .Y (n_4721));
  NAND4XL g175798(.A (n_2738), .B (n_2737), .C (n_2736), .D (n_3477),
       .Y (n_4720));
  NAND4XL g175799(.A (n_2702), .B (n_2701), .C (n_2700), .D (n_3476),
       .Y (n_4719));
  NAND4XL g175800(.A (n_2676), .B (n_2675), .C (n_2674), .D (n_3475),
       .Y (n_4718));
  NAND4XL g175801(.A (n_2637), .B (n_2636), .C (n_2635), .D (n_3474),
       .Y (n_4717));
  NAND4XL g175802(.A (n_2624), .B (n_2623), .C (n_2622), .D (n_3473),
       .Y (n_4716));
  OAI222X1 g175803(.A0 (n_762), .A1 (n_3236), .B0 (n_1802), .B1
       (n_3465), .C0 (n_683), .C1 (n_308), .Y (n_4715));
  OAI222X1 g175804(.A0 (n_583), .A1 (n_3236), .B0 (n_687), .B1
       (n_3465), .C0 (n_686), .C1 (n_308), .Y (n_4714));
  AOI222X1 g175805(.A0 (\cpuregs[2] [18]), .A1 (n_425), .B0
       (\cpuregs[15] [18]), .B1 (n_462), .C0 (\cpuregs[14] [18]), .C1
       (n_450), .Y (n_4713));
  MX2X1 g176402(.A (mem_do_rinst), .B (n_2613), .S0 (n_3396), .Y
       (n_4710));
  AOI221X1 g176403(.A0 (n_2615), .A1 (n_667), .B0 (instr_jalr), .B1
       (n_953), .C0 (n_3468), .Y (n_4709));
  OAI222X1 g176404(.A0 (n_611), .A1 (n_2151), .B0 (n_3248), .B1
       (n_2442), .C0 (n_651), .C1 (n_969), .Y (n_4708));
  OR4X1 g176405(.A (n_1346), .B (n_1354), .C (n_1348), .D (n_3169), .Y
       (n_4707));
  AOI22X1 g176406(.A0 (\cpuregs[16] [31]), .A1 (n_478), .B0
       (\cpuregs[17] [31]), .B1 (n_486), .Y (n_4706));
  AOI22X1 g176407(.A0 (\cpuregs[22] [31]), .A1 (n_482), .B0
       (\cpuregs[23] [31]), .B1 (n_464), .Y (n_4705));
  AOI22X1 g176408(.A0 (\cpuregs[20] [31]), .A1 (n_488), .B0
       (\cpuregs[21] [31]), .B1 (n_468), .Y (n_4704));
  AOI22X1 g176409(.A0 (\cpuregs[18] [31]), .A1 (n_492), .B0
       (\cpuregs[19] [31]), .B1 (n_502), .Y (n_4703));
  AOI22X1 g176410(.A0 (\cpuregs[24] [31]), .A1 (n_494), .B0
       (\cpuregs[25] [31]), .B1 (n_496), .Y (n_4702));
  AOI22X1 g176411(.A0 (\cpuregs[26] [31]), .A1 (n_490), .B0
       (\cpuregs[27] [31]), .B1 (n_498), .Y (n_4701));
  AOI22X1 g176412(.A0 (\cpuregs[28] [31]), .A1 (n_480), .B0
       (\cpuregs[29] [31]), .B1 (n_458), .Y (n_4700));
  AOI22X1 g176413(.A0 (\cpuregs[30] [31]), .A1 (n_500), .B0
       (\cpuregs[31] [31]), .B1 (n_476), .Y (n_4699));
  AOI22X1 g176414(.A0 (\cpuregs[8] [31]), .A1 (n_466), .B0
       (\cpuregs[12] [31]), .B1 (n_484), .Y (n_4698));
  AOI22X1 g176415(.A0 (\cpuregs[7] [31]), .A1 (n_474), .B0
       (\cpuregs[11] [31]), .B1 (n_448), .Y (n_4697));
  AOI22X1 g176416(.A0 (\cpuregs[9] [31]), .A1 (n_470), .B0
       (\cpuregs[10] [31]), .B1 (n_452), .Y (n_4696));
  AOI22X1 g176417(.A0 (\cpuregs[13] [31]), .A1 (n_454), .B0
       (\cpuregs[14] [31]), .B1 (n_450), .Y (n_4695));
  AOI22X1 g176418(.A0 (\cpuregs[2] [31]), .A1 (n_425), .B0
       (\cpuregs[15] [31]), .B1 (n_462), .Y (n_4694));
  AO22X1 g176419(.A0 (\cpuregs[5] [31]), .A1 (n_291), .B0
       (\cpuregs[6] [31]), .B1 (n_333), .Y (n_4693));
  AOI22X1 g176420(.A0 (\cpuregs[16] [30]), .A1 (n_478), .B0
       (\cpuregs[17] [30]), .B1 (n_486), .Y (n_4692));
  AOI22X1 g176421(.A0 (\cpuregs[22] [30]), .A1 (n_482), .B0
       (\cpuregs[23] [30]), .B1 (n_464), .Y (n_4691));
  AOI22X1 g176422(.A0 (\cpuregs[20] [30]), .A1 (n_488), .B0
       (\cpuregs[21] [30]), .B1 (n_468), .Y (n_4690));
  AOI22X1 g176423(.A0 (\cpuregs[18] [30]), .A1 (n_492), .B0
       (\cpuregs[19] [30]), .B1 (n_502), .Y (n_4689));
  AOI22X1 g176424(.A0 (\cpuregs[24] [30]), .A1 (n_494), .B0
       (\cpuregs[25] [30]), .B1 (n_496), .Y (n_4688));
  AOI22X1 g176425(.A0 (\cpuregs[30] [30]), .A1 (n_500), .B0
       (\cpuregs[31] [30]), .B1 (n_476), .Y (n_4687));
  AOI22X1 g176426(.A0 (\cpuregs[28] [30]), .A1 (n_480), .B0
       (\cpuregs[29] [30]), .B1 (n_458), .Y (n_4686));
  AOI22X1 g176427(.A0 (\cpuregs[26] [30]), .A1 (n_490), .B0
       (\cpuregs[27] [30]), .B1 (n_498), .Y (n_4685));
  AOI22X1 g176428(.A0 (\cpuregs[8] [30]), .A1 (n_466), .B0
       (\cpuregs[7] [30]), .B1 (n_474), .Y (n_4684));
  AOI22X1 g176429(.A0 (\cpuregs[9] [30]), .A1 (n_470), .B0
       (\cpuregs[10] [30]), .B1 (n_452), .Y (n_4683));
  AO22X1 g176430(.A0 (\cpuregs[11] [30]), .A1 (n_448), .B0
       (\cpuregs[14] [30]), .B1 (n_450), .Y (n_4682));
  AOI22X1 g176431(.A0 (\cpuregs[3] [30]), .A1 (n_423), .B0
       (\cpuregs[6] [30]), .B1 (n_333), .Y (n_4681));
  AOI22X1 g176432(.A0 (\cpuregs[4] [30]), .A1 (n_424), .B0
       (\cpuregs[5] [30]), .B1 (n_291), .Y (n_4680));
  AOI22X1 g176433(.A0 (\cpuregs[2] [30]), .A1 (n_425), .B0
       (\cpuregs[15] [30]), .B1 (n_462), .Y (n_4679));
  AOI22X1 g176434(.A0 (\cpuregs[16] [29]), .A1 (n_478), .B0
       (\cpuregs[17] [29]), .B1 (n_486), .Y (n_4678));
  AOI22X1 g176435(.A0 (\cpuregs[22] [29]), .A1 (n_482), .B0
       (\cpuregs[23] [29]), .B1 (n_464), .Y (n_4677));
  AOI22X1 g176436(.A0 (\cpuregs[20] [29]), .A1 (n_488), .B0
       (\cpuregs[21] [29]), .B1 (n_468), .Y (n_4676));
  AOI22X1 g176437(.A0 (\cpuregs[18] [29]), .A1 (n_492), .B0
       (\cpuregs[19] [29]), .B1 (n_502), .Y (n_4675));
  AOI22X1 g176438(.A0 (\cpuregs[26] [29]), .A1 (n_490), .B0
       (\cpuregs[31] [29]), .B1 (n_476), .Y (n_4674));
  AOI22X1 g176439(.A0 (\cpuregs[25] [29]), .A1 (n_496), .B0
       (\cpuregs[28] [29]), .B1 (n_480), .Y (n_4673));
  AOI22X1 g176440(.A0 (\cpuregs[29] [29]), .A1 (n_458), .B0
       (\cpuregs[30] [29]), .B1 (n_500), .Y (n_4672));
  AOI22X1 g176441(.A0 (\cpuregs[4] [29]), .A1 (n_424), .B0
       (\cpuregs[5] [29]), .B1 (n_291), .Y (n_4671));
  AOI22X1 g176442(.A0 (\cpuregs[12] [29]), .A1 (n_484), .B0
       (\cpuregs[13] [29]), .B1 (n_454), .Y (n_4670));
  AOI22X1 g176443(.A0 (\cpuregs[11] [29]), .A1 (n_448), .B0
       (\cpuregs[14] [29]), .B1 (n_450), .Y (n_4669));
  AO22X1 g176444(.A0 (\cpuregs[9] [29]), .A1 (n_470), .B0
       (\cpuregs[10] [29]), .B1 (n_452), .Y (n_4668));
  AOI22X1 g176445(.A0 (\cpuregs[24] [28]), .A1 (n_494), .B0
       (\cpuregs[25] [28]), .B1 (n_496), .Y (n_4667));
  AOI22X1 g176446(.A0 (\cpuregs[26] [28]), .A1 (n_490), .B0
       (\cpuregs[27] [28]), .B1 (n_498), .Y (n_4666));
  AOI22X1 g176447(.A0 (\cpuregs[28] [28]), .A1 (n_480), .B0
       (\cpuregs[29] [28]), .B1 (n_458), .Y (n_4665));
  AOI22X1 g176448(.A0 (\cpuregs[30] [28]), .A1 (n_500), .B0
       (\cpuregs[31] [28]), .B1 (n_476), .Y (n_4664));
  AOI22X1 g176449(.A0 (\cpuregs[20] [28]), .A1 (n_488), .B0
       (\cpuregs[19] [28]), .B1 (n_502), .Y (n_4663));
  AOI22X1 g176450(.A0 (\cpuregs[17] [28]), .A1 (n_486), .B0
       (\cpuregs[18] [28]), .B1 (n_492), .Y (n_4662));
  AOI22X1 g176451(.A0 (\cpuregs[16] [28]), .A1 (n_478), .B0
       (\cpuregs[23] [28]), .B1 (n_464), .Y (n_4661));
  AOI22X1 g176452(.A0 (\cpuregs[4] [28]), .A1 (n_424), .B0
       (\cpuregs[6] [28]), .B1 (n_333), .Y (n_4660));
  AO22X1 g176453(.A0 (\cpuregs[10] [28]), .A1 (n_452), .B0
       (\cpuregs[11] [28]), .B1 (n_448), .Y (n_4659));
  AOI22X1 g176454(.A0 (\cpuregs[8] [28]), .A1 (n_466), .B0
       (\cpuregs[7] [28]), .B1 (n_474), .Y (n_4658));
  AOI22X1 g176455(.A0 (\cpuregs[13] [28]), .A1 (n_454), .B0
       (\cpuregs[14] [28]), .B1 (n_450), .Y (n_4657));
  AOI22X1 g176456(.A0 (\cpuregs[16] [27]), .A1 (n_478), .B0
       (\cpuregs[17] [27]), .B1 (n_486), .Y (n_4656));
  AOI22X1 g176457(.A0 (\cpuregs[22] [27]), .A1 (n_482), .B0
       (\cpuregs[23] [27]), .B1 (n_464), .Y (n_4655));
  AOI22X1 g176458(.A0 (\cpuregs[20] [27]), .A1 (n_488), .B0
       (\cpuregs[21] [27]), .B1 (n_468), .Y (n_4654));
  AOI22X1 g176459(.A0 (\cpuregs[18] [27]), .A1 (n_492), .B0
       (\cpuregs[19] [27]), .B1 (n_502), .Y (n_4653));
  AOI22X1 g176460(.A0 (\cpuregs[25] [27]), .A1 (n_496), .B0
       (\cpuregs[28] [27]), .B1 (n_480), .Y (n_4652));
  AOI22X1 g176461(.A0 (\cpuregs[24] [27]), .A1 (n_494), .B0
       (\cpuregs[31] [27]), .B1 (n_476), .Y (n_4651));
  AOI22X1 g176462(.A0 (\cpuregs[27] [27]), .A1 (n_498), .B0
       (\cpuregs[30] [27]), .B1 (n_500), .Y (n_4650));
  AOI22X1 g176463(.A0 (\cpuregs[3] [27]), .A1 (n_423), .B0
       (\cpuregs[6] [27]), .B1 (n_333), .Y (n_4649));
  AO22X1 g176464(.A0 (\cpuregs[11] [27]), .A1 (n_448), .B0
       (\cpuregs[14] [27]), .B1 (n_450), .Y (n_4648));
  AOI22X1 g176465(.A0 (\cpuregs[8] [27]), .A1 (n_466), .B0
       (\cpuregs[7] [27]), .B1 (n_474), .Y (n_4647));
  AOI22X1 g176466(.A0 (\cpuregs[9] [27]), .A1 (n_470), .B0
       (\cpuregs[10] [27]), .B1 (n_452), .Y (n_4646));
  AOI22X1 g176467(.A0 (\cpuregs[16] [26]), .A1 (n_478), .B0
       (\cpuregs[17] [26]), .B1 (n_486), .Y (n_4645));
  AOI22X1 g176468(.A0 (\cpuregs[20] [26]), .A1 (n_488), .B0
       (\cpuregs[21] [26]), .B1 (n_468), .Y (n_4644));
  AOI22X1 g176469(.A0 (\cpuregs[18] [26]), .A1 (n_492), .B0
       (\cpuregs[19] [26]), .B1 (n_502), .Y (n_4643));
  AOI22X1 g176470(.A0 (\cpuregs[22] [26]), .A1 (n_482), .B0
       (\cpuregs[23] [26]), .B1 (n_464), .Y (n_4642));
  AOI22X1 g176471(.A0 (\cpuregs[25] [26]), .A1 (n_496), .B0
       (\cpuregs[28] [26]), .B1 (n_480), .Y (n_4641));
  AOI22X1 g176472(.A0 (\cpuregs[24] [26]), .A1 (n_494), .B0
       (\cpuregs[31] [26]), .B1 (n_476), .Y (n_4640));
  AOI22X1 g176473(.A0 (\cpuregs[27] [26]), .A1 (n_498), .B0
       (\cpuregs[30] [26]), .B1 (n_500), .Y (n_4639));
  AOI22X1 g176474(.A0 (\cpuregs[4] [26]), .A1 (n_424), .B0
       (\cpuregs[5] [26]), .B1 (n_291), .Y (n_4638));
  AO22X1 g176475(.A0 (\cpuregs[11] [26]), .A1 (n_448), .B0
       (\cpuregs[14] [26]), .B1 (n_450), .Y (n_4637));
  AOI22X1 g176476(.A0 (\cpuregs[8] [26]), .A1 (n_466), .B0
       (\cpuregs[7] [26]), .B1 (n_474), .Y (n_4636));
  AOI22X1 g176477(.A0 (\cpuregs[9] [26]), .A1 (n_470), .B0
       (\cpuregs[10] [26]), .B1 (n_452), .Y (n_4635));
  AOI22X1 g176478(.A0 (\cpuregs[16] [25]), .A1 (n_478), .B0
       (\cpuregs[17] [25]), .B1 (n_486), .Y (n_4634));
  AOI22X1 g176479(.A0 (\cpuregs[18] [25]), .A1 (n_492), .B0
       (\cpuregs[19] [25]), .B1 (n_502), .Y (n_4633));
  AOI22X1 g176480(.A0 (\cpuregs[20] [25]), .A1 (n_488), .B0
       (\cpuregs[21] [25]), .B1 (n_468), .Y (n_4632));
  AOI22X1 g176481(.A0 (\cpuregs[22] [25]), .A1 (n_482), .B0
       (\cpuregs[23] [25]), .B1 (n_464), .Y (n_4631));
  AOI22X1 g176482(.A0 (\cpuregs[24] [25]), .A1 (n_494), .B0
       (\cpuregs[25] [25]), .B1 (n_496), .Y (n_4630));
  AOI22X1 g176483(.A0 (\cpuregs[28] [25]), .A1 (n_480), .B0
       (\cpuregs[29] [25]), .B1 (n_458), .Y (n_4629));
  AOI22X1 g176484(.A0 (\cpuregs[26] [25]), .A1 (n_490), .B0
       (\cpuregs[27] [25]), .B1 (n_498), .Y (n_4628));
  AOI22X1 g176485(.A0 (\cpuregs[30] [25]), .A1 (n_500), .B0
       (\cpuregs[31] [25]), .B1 (n_476), .Y (n_4627));
  AOI22X1 g176486(.A0 (\cpuregs[8] [25]), .A1 (n_466), .B0
       (\cpuregs[12] [25]), .B1 (n_484), .Y (n_4626));
  AOI22X1 g176487(.A0 (\cpuregs[7] [25]), .A1 (n_474), .B0
       (\cpuregs[11] [25]), .B1 (n_448), .Y (n_4625));
  AOI22X1 g176488(.A0 (\cpuregs[9] [25]), .A1 (n_470), .B0
       (\cpuregs[10] [25]), .B1 (n_452), .Y (n_4624));
  AOI22X1 g176489(.A0 (\cpuregs[13] [25]), .A1 (n_454), .B0
       (\cpuregs[14] [25]), .B1 (n_450), .Y (n_4623));
  AOI22X1 g176490(.A0 (\cpuregs[4] [25]), .A1 (n_424), .B0
       (\cpuregs[3] [25]), .B1 (n_423), .Y (n_4622));
  AOI22X1 g176491(.A0 (\cpuregs[1] [25]), .A1 (n_456), .B0
       (\cpuregs[6] [25]), .B1 (n_333), .Y (n_4621));
  AOI22X1 g176492(.A0 (\cpuregs[16] [24]), .A1 (n_478), .B0
       (\cpuregs[17] [24]), .B1 (n_486), .Y (n_4620));
  AOI22X1 g176493(.A0 (\cpuregs[22] [24]), .A1 (n_482), .B0
       (\cpuregs[23] [24]), .B1 (n_464), .Y (n_4619));
  AOI22X1 g176494(.A0 (\cpuregs[20] [24]), .A1 (n_488), .B0
       (\cpuregs[21] [24]), .B1 (n_468), .Y (n_4618));
  AOI22X1 g176495(.A0 (\cpuregs[18] [24]), .A1 (n_492), .B0
       (\cpuregs[19] [24]), .B1 (n_502), .Y (n_4617));
  AOI22X1 g176496(.A0 (\cpuregs[29] [24]), .A1 (n_458), .B0
       (\cpuregs[30] [24]), .B1 (n_500), .Y (n_4616));
  AOI22X1 g176497(.A0 (\cpuregs[24] [24]), .A1 (n_494), .B0
       (\cpuregs[27] [24]), .B1 (n_498), .Y (n_4615));
  AOI22X1 g176498(.A0 (\cpuregs[25] [24]), .A1 (n_496), .B0
       (\cpuregs[28] [24]), .B1 (n_480), .Y (n_4614));
  AOI22X1 g176499(.A0 (\cpuregs[8] [24]), .A1 (n_466), .B0
       (\cpuregs[9] [24]), .B1 (n_470), .Y (n_4613));
  AOI22X1 g176500(.A0 (\cpuregs[10] [24]), .A1 (n_452), .B0
       (\cpuregs[7] [24]), .B1 (n_474), .Y (n_4612));
  AOI22X1 g176501(.A0 (\cpuregs[12] [24]), .A1 (n_484), .B0
       (\cpuregs[11] [24]), .B1 (n_448), .Y (n_4611));
  AOI22X1 g176502(.A0 (\cpuregs[13] [24]), .A1 (n_454), .B0
       (\cpuregs[14] [24]), .B1 (n_450), .Y (n_4610));
  AOI22X1 g176503(.A0 (\cpuregs[4] [24]), .A1 (n_424), .B0
       (\cpuregs[6] [24]), .B1 (n_333), .Y (n_4609));
  AOI22X1 g176504(.A0 (\cpuregs[1] [24]), .A1 (n_456), .B0
       (\cpuregs[2] [24]), .B1 (n_425), .Y (n_4608));
  AOI22X1 g176505(.A0 (\cpuregs[3] [24]), .A1 (n_423), .B0
       (\cpuregs[15] [24]), .B1 (n_462), .Y (n_4607));
  AOI22X1 g176506(.A0 (\cpuregs[24] [23]), .A1 (n_494), .B0
       (\cpuregs[25] [23]), .B1 (n_496), .Y (n_4606));
  AOI22X1 g176507(.A0 (\cpuregs[30] [23]), .A1 (n_500), .B0
       (\cpuregs[31] [23]), .B1 (n_476), .Y (n_4605));
  AO22X1 g176508(.A0 (\cpuregs[28] [23]), .A1 (n_480), .B0
       (\cpuregs[29] [23]), .B1 (n_458), .Y (n_4604));
  AOI22X1 g176509(.A0 (\cpuregs[18] [23]), .A1 (n_492), .B0
       (\cpuregs[19] [23]), .B1 (n_502), .Y (n_4603));
  AOI22X1 g176510(.A0 (\cpuregs[16] [23]), .A1 (n_478), .B0
       (\cpuregs[17] [23]), .B1 (n_486), .Y (n_4602));
  AOI22X1 g176511(.A0 (\cpuregs[20] [23]), .A1 (n_488), .B0
       (\cpuregs[21] [23]), .B1 (n_468), .Y (n_4601));
  AOI22X1 g176512(.A0 (\cpuregs[8] [23]), .A1 (n_466), .B0
       (\cpuregs[7] [23]), .B1 (n_474), .Y (n_4600));
  AOI22X1 g176513(.A0 (\cpuregs[12] [23]), .A1 (n_484), .B0
       (\cpuregs[11] [23]), .B1 (n_448), .Y (n_4599));
  AOI22X1 g176514(.A0 (\cpuregs[9] [23]), .A1 (n_470), .B0
       (\cpuregs[13] [23]), .B1 (n_454), .Y (n_4598));
  AOI22X1 g176515(.A0 (\cpuregs[10] [23]), .A1 (n_452), .B0
       (\cpuregs[14] [23]), .B1 (n_450), .Y (n_4597));
  AOI22X1 g176516(.A0 (\cpuregs[18] [22]), .A1 (n_492), .B0
       (\cpuregs[19] [22]), .B1 (n_502), .Y (n_4596));
  AOI22X1 g176517(.A0 (\cpuregs[16] [22]), .A1 (n_478), .B0
       (\cpuregs[17] [22]), .B1 (n_486), .Y (n_4595));
  AOI22X1 g176518(.A0 (\cpuregs[20] [22]), .A1 (n_488), .B0
       (\cpuregs[21] [22]), .B1 (n_468), .Y (n_4594));
  AOI22X1 g176519(.A0 (\cpuregs[22] [22]), .A1 (n_482), .B0
       (\cpuregs[23] [22]), .B1 (n_464), .Y (n_4593));
  AOI22X1 g176520(.A0 (\cpuregs[9] [22]), .A1 (n_470), .B0
       (\cpuregs[12] [22]), .B1 (n_484), .Y (n_4592));
  AOI22X1 g176521(.A0 (\cpuregs[10] [22]), .A1 (n_452), .B0
       (\cpuregs[11] [22]), .B1 (n_448), .Y (n_4591));
  AOI22X1 g176522(.A0 (\cpuregs[13] [22]), .A1 (n_454), .B0
       (\cpuregs[14] [22]), .B1 (n_450), .Y (n_4590));
  AOI22X1 g176523(.A0 (\cpuregs[24] [22]), .A1 (n_494), .B0
       (\cpuregs[25] [22]), .B1 (n_496), .Y (n_4589));
  AOI22X1 g176524(.A0 (\cpuregs[30] [22]), .A1 (n_500), .B0
       (\cpuregs[31] [22]), .B1 (n_476), .Y (n_4588));
  AOI22X1 g176525(.A0 (\cpuregs[28] [22]), .A1 (n_480), .B0
       (\cpuregs[29] [22]), .B1 (n_458), .Y (n_4587));
  AOI22X1 g176526(.A0 (\cpuregs[26] [22]), .A1 (n_490), .B0
       (\cpuregs[27] [22]), .B1 (n_498), .Y (n_4586));
  AOI22X1 g176527(.A0 (\cpuregs[16] [21]), .A1 (n_478), .B0
       (\cpuregs[17] [21]), .B1 (n_486), .Y (n_4585));
  AOI22X1 g176528(.A0 (\cpuregs[18] [21]), .A1 (n_492), .B0
       (\cpuregs[19] [21]), .B1 (n_502), .Y (n_4584));
  AOI22X1 g176529(.A0 (\cpuregs[20] [21]), .A1 (n_488), .B0
       (\cpuregs[21] [21]), .B1 (n_468), .Y (n_4583));
  AOI22X1 g176530(.A0 (\cpuregs[22] [21]), .A1 (n_482), .B0
       (\cpuregs[23] [21]), .B1 (n_464), .Y (n_4582));
  AOI22X1 g176531(.A0 (\cpuregs[24] [21]), .A1 (n_494), .B0
       (\cpuregs[25] [21]), .B1 (n_496), .Y (n_4581));
  AOI22X1 g176532(.A0 (\cpuregs[28] [21]), .A1 (n_480), .B0
       (\cpuregs[29] [21]), .B1 (n_458), .Y (n_4580));
  AOI22X1 g176533(.A0 (\cpuregs[26] [21]), .A1 (n_490), .B0
       (\cpuregs[27] [21]), .B1 (n_498), .Y (n_4579));
  AOI22X1 g176534(.A0 (\cpuregs[30] [21]), .A1 (n_500), .B0
       (\cpuregs[31] [21]), .B1 (n_476), .Y (n_4578));
  AO22X1 g176535(.A0 (\cpuregs[10] [21]), .A1 (n_452), .B0
       (\cpuregs[13] [21]), .B1 (n_454), .Y (n_4577));
  AOI22X1 g176536(.A0 (\cpuregs[8] [21]), .A1 (n_466), .B0
       (\cpuregs[11] [21]), .B1 (n_448), .Y (n_4576));
  AOI22X1 g176537(.A0 (\cpuregs[12] [21]), .A1 (n_484), .B0
       (\cpuregs[14] [21]), .B1 (n_450), .Y (n_4575));
  AOI22X1 g176538(.A0 (\cpuregs[16] [20]), .A1 (n_478), .B0
       (\cpuregs[17] [20]), .B1 (n_486), .Y (n_4574));
  AOI22X1 g176539(.A0 (\cpuregs[22] [20]), .A1 (n_482), .B0
       (\cpuregs[23] [20]), .B1 (n_464), .Y (n_4573));
  AOI22X1 g176540(.A0 (\cpuregs[20] [20]), .A1 (n_488), .B0
       (\cpuregs[21] [20]), .B1 (n_468), .Y (n_4572));
  AOI22X1 g176541(.A0 (\cpuregs[18] [20]), .A1 (n_492), .B0
       (\cpuregs[19] [20]), .B1 (n_502), .Y (n_4571));
  AOI22X1 g176542(.A0 (\cpuregs[24] [20]), .A1 (n_494), .B0
       (\cpuregs[25] [20]), .B1 (n_496), .Y (n_4570));
  AOI22X1 g176543(.A0 (\cpuregs[28] [20]), .A1 (n_480), .B0
       (\cpuregs[29] [20]), .B1 (n_458), .Y (n_4569));
  AOI22X1 g176544(.A0 (\cpuregs[26] [20]), .A1 (n_490), .B0
       (\cpuregs[27] [20]), .B1 (n_498), .Y (n_4568));
  AOI22X1 g176545(.A0 (\cpuregs[30] [20]), .A1 (n_500), .B0
       (\cpuregs[31] [20]), .B1 (n_476), .Y (n_4567));
  AOI22X1 g176546(.A0 (\cpuregs[8] [20]), .A1 (n_466), .B0
       (\cpuregs[7] [20]), .B1 (n_474), .Y (n_4566));
  AOI22X1 g176547(.A0 (\cpuregs[12] [20]), .A1 (n_484), .B0
       (\cpuregs[11] [20]), .B1 (n_448), .Y (n_4565));
  AOI22X1 g176548(.A0 (\cpuregs[9] [20]), .A1 (n_470), .B0
       (\cpuregs[13] [20]), .B1 (n_454), .Y (n_4564));
  AOI22X1 g176549(.A0 (\cpuregs[10] [20]), .A1 (n_452), .B0
       (\cpuregs[14] [20]), .B1 (n_450), .Y (n_4563));
  AOI22X1 g176550(.A0 (\cpuregs[4] [20]), .A1 (n_424), .B0
       (\cpuregs[6] [20]), .B1 (n_333), .Y (n_4562));
  AOI22X1 g176551(.A0 (\cpuregs[2] [20]), .A1 (n_425), .B0
       (\cpuregs[3] [20]), .B1 (n_423), .Y (n_4561));
  AOI22X1 g176552(.A0 (\cpuregs[24] [19]), .A1 (n_494), .B0
       (\cpuregs[25] [19]), .B1 (n_496), .Y (n_4560));
  AOI22X1 g176553(.A0 (\cpuregs[30] [19]), .A1 (n_500), .B0
       (\cpuregs[31] [19]), .B1 (n_476), .Y (n_4559));
  AOI22X1 g176554(.A0 (\cpuregs[28] [19]), .A1 (n_480), .B0
       (\cpuregs[29] [19]), .B1 (n_458), .Y (n_4558));
  AOI22X1 g176555(.A0 (\cpuregs[26] [19]), .A1 (n_490), .B0
       (\cpuregs[27] [19]), .B1 (n_498), .Y (n_4557));
  AOI22X1 g176556(.A0 (\cpuregs[18] [19]), .A1 (n_492), .B0
       (\cpuregs[19] [19]), .B1 (n_502), .Y (n_4556));
  AOI22X1 g176557(.A0 (\cpuregs[16] [19]), .A1 (n_478), .B0
       (\cpuregs[17] [19]), .B1 (n_486), .Y (n_4555));
  AOI22X1 g176558(.A0 (\cpuregs[22] [19]), .A1 (n_482), .B0
       (\cpuregs[23] [19]), .B1 (n_464), .Y (n_4554));
  AOI22X1 g176559(.A0 (\cpuregs[9] [19]), .A1 (n_470), .B0
       (\cpuregs[10] [19]), .B1 (n_452), .Y (n_4553));
  AOI22X1 g176560(.A0 (\cpuregs[12] [19]), .A1 (n_484), .B0
       (\cpuregs[11] [19]), .B1 (n_448), .Y (n_4552));
  AOI22X1 g176561(.A0 (\cpuregs[8] [19]), .A1 (n_466), .B0
       (\cpuregs[13] [19]), .B1 (n_454), .Y (n_4551));
  AOI22X1 g176562(.A0 (\cpuregs[7] [19]), .A1 (n_474), .B0
       (\cpuregs[14] [19]), .B1 (n_450), .Y (n_4550));
  AOI22X1 g176563(.A0 (\cpuregs[1] [18]), .A1 (n_456), .B0
       (\cpuregs[8] [18]), .B1 (n_466), .Y (n_4549));
  AOI22X1 g176564(.A0 (\cpuregs[12] [18]), .A1 (n_484), .B0
       (\cpuregs[11] [18]), .B1 (n_448), .Y (n_4548));
  AO22X1 g176565(.A0 (\cpuregs[10] [18]), .A1 (n_452), .B0
       (\cpuregs[13] [18]), .B1 (n_454), .Y (n_4547));
  AOI22X1 g176566(.A0 (\cpuregs[16] [18]), .A1 (n_478), .B0
       (\cpuregs[17] [18]), .B1 (n_486), .Y (n_4546));
  AOI22X1 g176567(.A0 (\cpuregs[18] [18]), .A1 (n_492), .B0
       (\cpuregs[19] [18]), .B1 (n_502), .Y (n_4545));
  AOI22X1 g176568(.A0 (\cpuregs[20] [18]), .A1 (n_488), .B0
       (\cpuregs[21] [18]), .B1 (n_468), .Y (n_4544));
  AOI22X1 g176569(.A0 (\cpuregs[22] [18]), .A1 (n_482), .B0
       (\cpuregs[23] [18]), .B1 (n_464), .Y (n_4543));
  AOI22X1 g176570(.A0 (\cpuregs[5] [18]), .A1 (n_291), .B0
       (\cpuregs[6] [18]), .B1 (n_333), .Y (n_4542));
  AOI22X1 g176571(.A0 (\cpuregs[3] [18]), .A1 (n_423), .B0 (n_833), .B1
       (n_50), .Y (n_4541));
  AOI22X1 g176572(.A0 (\cpuregs[24] [18]), .A1 (n_494), .B0
       (\cpuregs[25] [18]), .B1 (n_496), .Y (n_4540));
  AOI22X1 g176573(.A0 (\cpuregs[26] [18]), .A1 (n_490), .B0
       (\cpuregs[27] [18]), .B1 (n_498), .Y (n_4539));
  AOI22X1 g176574(.A0 (\cpuregs[30] [18]), .A1 (n_500), .B0
       (\cpuregs[31] [18]), .B1 (n_476), .Y (n_4538));
  AOI22X1 g176575(.A0 (\cpuregs[28] [18]), .A1 (n_480), .B0
       (\cpuregs[29] [18]), .B1 (n_458), .Y (n_4537));
  AOI22X1 g176576(.A0 (\cpuregs[16] [17]), .A1 (n_478), .B0
       (\cpuregs[17] [17]), .B1 (n_486), .Y (n_4536));
  NAND2X1 g176577(.A (n_2441), .B (n_310), .Y (n_4535));
  NAND2X1 g176578(.A (n_0), .B (n_4288), .Y (n_4534));
  NAND2X1 g176579(.A (n_326), .B (n_4289), .Y (n_4533));
  OAI221X1 g176580(.A0 (n_683), .A1 (n_3253), .B0 (n_593), .B1 (n_667),
       .C0 (n_2170), .Y (n_4532));
  AOI22X1 g176581(.A0 (\cpuregs[18] [17]), .A1 (n_492), .B0
       (\cpuregs[19] [17]), .B1 (n_502), .Y (n_4531));
  NOR4X1 g176582(.A (\reg_op2[8]_9677 ), .B (\reg_op2[13]_9682 ), .C
       (\reg_op2[14]_9683 ), .D (n_3171), .Y (n_4530));
  NAND4XL g176583(.A (n_1356), .B (n_1323), .C (n_323), .D (n_3251), .Y
       (n_4529));
  OAI2BB1X1 g176584(.A0N (decoded_imm[2]), .A1N (n_421), .B0 (n_4085),
       .Y (n_4528));
  OAI2BB1X1 g176585(.A0N (decoded_imm[3]), .A1N (n_421), .B0 (n_4084),
       .Y (n_4527));
  AOI211XL g176586(.A0 (\cpuregs[3] [7]), .A1 (n_2503), .B0 (n_3256),
       .C0 (n_3124), .Y (n_4526));
  AOI211XL g176587(.A0 (\cpuregs[5] [24]), .A1 (n_2492), .B0 (n_3255),
       .C0 (n_3091), .Y (n_4525));
  AOI211XL g176588(.A0 (\cpuregs[3] [29]), .A1 (n_2503), .B0 (n_3395),
       .C0 (n_3131), .Y (n_4524));
  AOI22X1 g176589(.A0 (\cpuregs[9] [0]), .A1 (n_470), .B0
       (\cpuregs[10] [0]), .B1 (n_452), .Y (n_4523));
  AOI22X1 g176590(.A0 (\cpuregs[8] [0]), .A1 (n_466), .B0
       (\cpuregs[7] [0]), .B1 (n_474), .Y (n_4522));
  AO22X1 g176591(.A0 (\cpuregs[11] [0]), .A1 (n_448), .B0
       (\cpuregs[14] [0]), .B1 (n_450), .Y (n_4521));
  AOI22X1 g176592(.A0 (\cpuregs[3] [0]), .A1 (n_423), .B0
       (\cpuregs[6] [0]), .B1 (n_333), .Y (n_4520));
  AOI22X1 g176593(.A0 (\cpuregs[20] [0]), .A1 (n_488), .B0
       (\cpuregs[23] [0]), .B1 (n_464), .Y (n_4519));
  AOI22X1 g176594(.A0 (\cpuregs[18] [0]), .A1 (n_492), .B0
       (\cpuregs[21] [0]), .B1 (n_468), .Y (n_4518));
  AOI22X1 g176595(.A0 (\cpuregs[16] [0]), .A1 (n_478), .B0
       (\cpuregs[19] [0]), .B1 (n_502), .Y (n_4517));
  AOI22X1 g176596(.A0 (\cpuregs[30] [0]), .A1 (n_500), .B0
       (\cpuregs[31] [0]), .B1 (n_476), .Y (n_4516));
  AOI22X1 g176597(.A0 (\cpuregs[28] [0]), .A1 (n_480), .B0
       (\cpuregs[29] [0]), .B1 (n_458), .Y (n_4515));
  AOI22X1 g176598(.A0 (\cpuregs[26] [0]), .A1 (n_490), .B0
       (\cpuregs[27] [0]), .B1 (n_498), .Y (n_4514));
  AOI22X1 g176599(.A0 (\cpuregs[24] [0]), .A1 (n_494), .B0
       (\cpuregs[25] [0]), .B1 (n_496), .Y (n_4513));
  AOI22X1 g176600(.A0 (\cpuregs[26] [1]), .A1 (n_490), .B0
       (\cpuregs[27] [1]), .B1 (n_498), .Y (n_4512));
  AOI22X1 g176601(.A0 (\cpuregs[24] [1]), .A1 (n_494), .B0
       (\cpuregs[25] [1]), .B1 (n_496), .Y (n_4511));
  AOI22X1 g176602(.A0 (\cpuregs[28] [1]), .A1 (n_480), .B0
       (\cpuregs[29] [1]), .B1 (n_458), .Y (n_4510));
  AOI22X1 g176603(.A0 (\cpuregs[18] [1]), .A1 (n_492), .B0
       (\cpuregs[19] [1]), .B1 (n_502), .Y (n_4509));
  AOI22X1 g176604(.A0 (\cpuregs[20] [1]), .A1 (n_488), .B0
       (\cpuregs[21] [1]), .B1 (n_468), .Y (n_4508));
  AOI22X1 g176605(.A0 (\cpuregs[22] [1]), .A1 (n_482), .B0
       (\cpuregs[23] [1]), .B1 (n_464), .Y (n_4507));
  AOI22X1 g176606(.A0 (\cpuregs[16] [1]), .A1 (n_478), .B0
       (\cpuregs[17] [1]), .B1 (n_486), .Y (n_4506));
  AOI22X1 g176607(.A0 (\cpuregs[15] [1]), .A1 (n_462), .B0 (n_833), .B1
       (n_62), .Y (n_4505));
  AOI22X1 g176608(.A0 (\cpuregs[3] [1]), .A1 (n_423), .B0
       (\cpuregs[6] [1]), .B1 (n_333), .Y (n_4504));
  AOI22X1 g176609(.A0 (\cpuregs[1] [1]), .A1 (n_456), .B0 (reg_pc[1]),
       .B1 (n_961), .Y (n_4503));
  AOI22X1 g176610(.A0 (\cpuregs[13] [1]), .A1 (n_454), .B0
       (\cpuregs[14] [1]), .B1 (n_450), .Y (n_4502));
  AOI22X1 g176611(.A0 (\cpuregs[12] [1]), .A1 (n_484), .B0
       (\cpuregs[11] [1]), .B1 (n_448), .Y (n_4501));
  AOI22X1 g176612(.A0 (\cpuregs[10] [1]), .A1 (n_452), .B0
       (\cpuregs[7] [1]), .B1 (n_474), .Y (n_4500));
  AOI22X1 g176613(.A0 (\cpuregs[8] [1]), .A1 (n_466), .B0
       (\cpuregs[9] [1]), .B1 (n_470), .Y (n_4499));
  AO22X1 g176614(.A0 (\cpuregs[5] [2]), .A1 (n_291), .B0
       (\cpuregs[6] [2]), .B1 (n_333), .Y (n_4498));
  AOI22X1 g176615(.A0 (\cpuregs[2] [2]), .A1 (n_425), .B0
       (\cpuregs[15] [2]), .B1 (n_462), .Y (n_4497));
  AOI22X1 g176616(.A0 (\cpuregs[30] [2]), .A1 (n_500), .B0
       (\cpuregs[31] [2]), .B1 (n_476), .Y (n_4496));
  AOI22X1 g176617(.A0 (\cpuregs[28] [2]), .A1 (n_480), .B0
       (\cpuregs[29] [2]), .B1 (n_458), .Y (n_4495));
  AOI22X1 g176618(.A0 (\cpuregs[26] [2]), .A1 (n_490), .B0
       (\cpuregs[27] [2]), .B1 (n_498), .Y (n_4494));
  AOI22X1 g176619(.A0 (\cpuregs[24] [2]), .A1 (n_494), .B0
       (\cpuregs[25] [2]), .B1 (n_496), .Y (n_4493));
  AOI22X1 g176620(.A0 (\cpuregs[22] [2]), .A1 (n_482), .B0
       (\cpuregs[23] [2]), .B1 (n_464), .Y (n_4492));
  AOI22X1 g176621(.A0 (\cpuregs[18] [2]), .A1 (n_492), .B0
       (\cpuregs[19] [2]), .B1 (n_502), .Y (n_4491));
  AOI22X1 g176622(.A0 (\cpuregs[20] [2]), .A1 (n_488), .B0
       (\cpuregs[21] [2]), .B1 (n_468), .Y (n_4490));
  AOI22X1 g176623(.A0 (\cpuregs[16] [2]), .A1 (n_478), .B0
       (\cpuregs[17] [2]), .B1 (n_486), .Y (n_4489));
  AOI22X1 g176624(.A0 (\cpuregs[10] [2]), .A1 (n_452), .B0
       (\cpuregs[14] [2]), .B1 (n_450), .Y (n_4488));
  AOI22X1 g176625(.A0 (\cpuregs[9] [2]), .A1 (n_470), .B0
       (\cpuregs[13] [2]), .B1 (n_454), .Y (n_4487));
  AOI22X1 g176626(.A0 (\cpuregs[12] [2]), .A1 (n_484), .B0
       (\cpuregs[11] [2]), .B1 (n_448), .Y (n_4486));
  AOI22X1 g176627(.A0 (\cpuregs[8] [2]), .A1 (n_466), .B0
       (\cpuregs[7] [2]), .B1 (n_474), .Y (n_4485));
  AOI22X1 g176628(.A0 (\cpuregs[5] [3]), .A1 (n_291), .B0
       (\cpuregs[6] [3]), .B1 (n_333), .Y (n_4484));
  AOI22X1 g176629(.A0 (\cpuregs[4] [3]), .A1 (n_424), .B0
       (\cpuregs[3] [3]), .B1 (n_423), .Y (n_4483));
  AOI22X1 g176630(.A0 (\cpuregs[7] [3]), .A1 (n_474), .B0
       (\cpuregs[14] [3]), .B1 (n_450), .Y (n_4482));
  AOI22X1 g176631(.A0 (\cpuregs[8] [3]), .A1 (n_466), .B0
       (\cpuregs[13] [3]), .B1 (n_454), .Y (n_4481));
  AOI22X1 g176632(.A0 (\cpuregs[12] [3]), .A1 (n_484), .B0
       (\cpuregs[11] [3]), .B1 (n_448), .Y (n_4480));
  AOI22X1 g176633(.A0 (\cpuregs[9] [3]), .A1 (n_470), .B0
       (\cpuregs[10] [3]), .B1 (n_452), .Y (n_4479));
  AOI22X1 g176634(.A0 (\cpuregs[30] [3]), .A1 (n_500), .B0
       (\cpuregs[31] [3]), .B1 (n_476), .Y (n_4478));
  AOI22X1 g176635(.A0 (\cpuregs[26] [3]), .A1 (n_490), .B0
       (\cpuregs[27] [3]), .B1 (n_498), .Y (n_4477));
  AOI22X1 g176636(.A0 (\cpuregs[28] [3]), .A1 (n_480), .B0
       (\cpuregs[29] [3]), .B1 (n_458), .Y (n_4476));
  AOI22X1 g176637(.A0 (\cpuregs[24] [3]), .A1 (n_494), .B0
       (\cpuregs[25] [3]), .B1 (n_496), .Y (n_4475));
  AOI22X1 g176638(.A0 (\cpuregs[22] [3]), .A1 (n_482), .B0
       (\cpuregs[23] [3]), .B1 (n_464), .Y (n_4474));
  AOI22X1 g176639(.A0 (\cpuregs[20] [3]), .A1 (n_488), .B0
       (\cpuregs[21] [3]), .B1 (n_468), .Y (n_4473));
  AOI22X1 g176640(.A0 (\cpuregs[18] [3]), .A1 (n_492), .B0
       (\cpuregs[19] [3]), .B1 (n_502), .Y (n_4472));
  AOI22X1 g176641(.A0 (\cpuregs[16] [3]), .A1 (n_478), .B0
       (\cpuregs[17] [3]), .B1 (n_486), .Y (n_4471));
  AOI22X1 g176642(.A0 (\cpuregs[3] [4]), .A1 (n_423), .B0
       (\cpuregs[15] [4]), .B1 (n_462), .Y (n_4470));
  AOI22X1 g176643(.A0 (\cpuregs[1] [4]), .A1 (n_456), .B0
       (\cpuregs[2] [4]), .B1 (n_425), .Y (n_4469));
  AOI22X1 g176644(.A0 (\cpuregs[4] [4]), .A1 (n_424), .B0
       (\cpuregs[6] [4]), .B1 (n_333), .Y (n_4468));
  AOI22X1 g176645(.A0 (\cpuregs[7] [4]), .A1 (n_474), .B0
       (\cpuregs[14] [4]), .B1 (n_450), .Y (n_4467));
  AOI22X1 g176646(.A0 (\cpuregs[8] [4]), .A1 (n_466), .B0
       (\cpuregs[13] [4]), .B1 (n_454), .Y (n_4466));
  AOI22X1 g176647(.A0 (\cpuregs[12] [4]), .A1 (n_484), .B0
       (\cpuregs[11] [4]), .B1 (n_448), .Y (n_4465));
  AOI22X1 g176648(.A0 (\cpuregs[9] [4]), .A1 (n_470), .B0
       (\cpuregs[10] [4]), .B1 (n_452), .Y (n_4464));
  AOI22X1 g176649(.A0 (\cpuregs[27] [4]), .A1 (n_498), .B0
       (\cpuregs[30] [4]), .B1 (n_500), .Y (n_4463));
  AOI22X1 g176650(.A0 (\cpuregs[24] [4]), .A1 (n_494), .B0
       (\cpuregs[31] [4]), .B1 (n_476), .Y (n_4462));
  AOI22X1 g176651(.A0 (\cpuregs[25] [4]), .A1 (n_496), .B0
       (\cpuregs[28] [4]), .B1 (n_480), .Y (n_4461));
  AOI22X1 g176652(.A0 (\cpuregs[22] [4]), .A1 (n_482), .B0
       (\cpuregs[23] [4]), .B1 (n_464), .Y (n_4460));
  AOI22X1 g176653(.A0 (\cpuregs[18] [4]), .A1 (n_492), .B0
       (\cpuregs[19] [4]), .B1 (n_502), .Y (n_4459));
  AOI22X1 g176654(.A0 (\cpuregs[20] [4]), .A1 (n_488), .B0
       (\cpuregs[21] [4]), .B1 (n_468), .Y (n_4458));
  AOI22X1 g176655(.A0 (\cpuregs[16] [4]), .A1 (n_478), .B0
       (\cpuregs[17] [4]), .B1 (n_486), .Y (n_4457));
  AOI22X1 g176656(.A0 (\cpuregs[13] [5]), .A1 (n_454), .B0
       (\cpuregs[14] [5]), .B1 (n_450), .Y (n_4456));
  AOI22X1 g176657(.A0 (\cpuregs[12] [5]), .A1 (n_484), .B0
       (\cpuregs[11] [5]), .B1 (n_448), .Y (n_4455));
  AO22X1 g176658(.A0 (\cpuregs[8] [5]), .A1 (n_466), .B0
       (\cpuregs[9] [5]), .B1 (n_470), .Y (n_4454));
  AOI22X1 g176659(.A0 (\cpuregs[4] [5]), .A1 (n_424), .B0
       (\cpuregs[6] [5]), .B1 (n_333), .Y (n_4453));
  AOI22X1 g176660(.A0 (\cpuregs[19] [5]), .A1 (n_502), .B0
       (\cpuregs[22] [5]), .B1 (n_482), .Y (n_4452));
  AOI22X1 g176661(.A0 (\cpuregs[16] [5]), .A1 (n_478), .B0
       (\cpuregs[23] [5]), .B1 (n_464), .Y (n_4451));
  AOI22X1 g176662(.A0 (\cpuregs[17] [5]), .A1 (n_486), .B0
       (\cpuregs[20] [5]), .B1 (n_488), .Y (n_4450));
  AOI22X1 g176663(.A0 (\cpuregs[26] [5]), .A1 (n_490), .B0
       (\cpuregs[27] [5]), .B1 (n_498), .Y (n_4449));
  AOI22X1 g176664(.A0 (\cpuregs[28] [5]), .A1 (n_480), .B0
       (\cpuregs[29] [5]), .B1 (n_458), .Y (n_4448));
  AOI22X1 g176665(.A0 (\cpuregs[30] [5]), .A1 (n_500), .B0
       (\cpuregs[31] [5]), .B1 (n_476), .Y (n_4447));
  AOI22X1 g176666(.A0 (\cpuregs[24] [5]), .A1 (n_494), .B0
       (\cpuregs[25] [5]), .B1 (n_496), .Y (n_4446));
  AOI22X1 g176667(.A0 (\cpuregs[18] [6]), .A1 (n_492), .B0
       (\cpuregs[19] [6]), .B1 (n_502), .Y (n_4445));
  AOI22X1 g176668(.A0 (\cpuregs[20] [6]), .A1 (n_488), .B0
       (\cpuregs[21] [6]), .B1 (n_468), .Y (n_4444));
  AO22X1 g176669(.A0 (\cpuregs[16] [6]), .A1 (n_478), .B0
       (\cpuregs[17] [6]), .B1 (n_486), .Y (n_4443));
  AOI22X1 g176670(.A0 (\cpuregs[30] [6]), .A1 (n_500), .B0
       (\cpuregs[31] [6]), .B1 (n_476), .Y (n_4442));
  AOI22X1 g176671(.A0 (\cpuregs[28] [6]), .A1 (n_480), .B0
       (\cpuregs[29] [6]), .B1 (n_458), .Y (n_4441));
  AOI22X1 g176672(.A0 (\cpuregs[26] [6]), .A1 (n_490), .B0
       (\cpuregs[27] [6]), .B1 (n_498), .Y (n_4440));
  AOI22X1 g176673(.A0 (\cpuregs[24] [6]), .A1 (n_494), .B0
       (\cpuregs[25] [6]), .B1 (n_496), .Y (n_4439));
  AOI22X1 g176674(.A0 (\cpuregs[4] [6]), .A1 (n_424), .B0
       (\cpuregs[3] [6]), .B1 (n_423), .Y (n_4438));
  AOI22X1 g176675(.A0 (\cpuregs[5] [6]), .A1 (n_291), .B0
       (\cpuregs[6] [6]), .B1 (n_333), .Y (n_4437));
  AOI22X1 g176676(.A0 (\cpuregs[9] [6]), .A1 (n_470), .B0
       (\cpuregs[13] [6]), .B1 (n_454), .Y (n_4436));
  AOI22X1 g176677(.A0 (\cpuregs[10] [6]), .A1 (n_452), .B0
       (\cpuregs[14] [6]), .B1 (n_450), .Y (n_4435));
  AOI22X1 g176678(.A0 (\cpuregs[12] [6]), .A1 (n_484), .B0
       (\cpuregs[11] [6]), .B1 (n_448), .Y (n_4434));
  AOI22X1 g176679(.A0 (\cpuregs[8] [6]), .A1 (n_466), .B0
       (\cpuregs[7] [6]), .B1 (n_474), .Y (n_4433));
  AOI22X1 g176680(.A0 (\cpuregs[10] [7]), .A1 (n_452), .B0
       (\cpuregs[14] [7]), .B1 (n_450), .Y (n_4432));
  AOI22X1 g176681(.A0 (\cpuregs[9] [7]), .A1 (n_470), .B0
       (\cpuregs[13] [7]), .B1 (n_454), .Y (n_4431));
  AOI22X1 g176682(.A0 (\cpuregs[12] [7]), .A1 (n_484), .B0
       (\cpuregs[11] [7]), .B1 (n_448), .Y (n_4430));
  AOI22X1 g176683(.A0 (\cpuregs[8] [7]), .A1 (n_466), .B0
       (\cpuregs[7] [7]), .B1 (n_474), .Y (n_4429));
  AO22X1 g176684(.A0 (\cpuregs[20] [7]), .A1 (n_488), .B0
       (\cpuregs[21] [7]), .B1 (n_468), .Y (n_4428));
  AOI22X1 g176685(.A0 (\cpuregs[22] [7]), .A1 (n_482), .B0
       (\cpuregs[23] [7]), .B1 (n_464), .Y (n_4427));
  AOI22X1 g176686(.A0 (\cpuregs[30] [7]), .A1 (n_500), .B0
       (\cpuregs[31] [7]), .B1 (n_476), .Y (n_4426));
  AOI22X1 g176687(.A0 (\cpuregs[28] [7]), .A1 (n_480), .B0
       (\cpuregs[29] [7]), .B1 (n_458), .Y (n_4425));
  AOI22X1 g176688(.A0 (\cpuregs[26] [7]), .A1 (n_490), .B0
       (\cpuregs[27] [7]), .B1 (n_498), .Y (n_4424));
  AOI22X1 g176689(.A0 (\cpuregs[24] [7]), .A1 (n_494), .B0
       (\cpuregs[25] [7]), .B1 (n_496), .Y (n_4423));
  AOI22X1 g176690(.A0 (\cpuregs[3] [8]), .A1 (n_423), .B0
       (\cpuregs[15] [8]), .B1 (n_462), .Y (n_4422));
  AOI22X1 g176691(.A0 (\cpuregs[1] [8]), .A1 (n_456), .B0
       (\cpuregs[2] [8]), .B1 (n_425), .Y (n_4421));
  AOI22X1 g176692(.A0 (\cpuregs[4] [8]), .A1 (n_424), .B0
       (\cpuregs[6] [8]), .B1 (n_333), .Y (n_4420));
  AOI22X1 g176693(.A0 (\cpuregs[8] [8]), .A1 (n_466), .B0
       (\cpuregs[7] [8]), .B1 (n_474), .Y (n_4419));
  AOI22X1 g176694(.A0 (\cpuregs[13] [8]), .A1 (n_454), .B0
       (\cpuregs[14] [8]), .B1 (n_450), .Y (n_4418));
  AOI22X1 g176695(.A0 (\cpuregs[10] [8]), .A1 (n_452), .B0
       (\cpuregs[11] [8]), .B1 (n_448), .Y (n_4417));
  AOI22X1 g176696(.A0 (\cpuregs[9] [8]), .A1 (n_470), .B0
       (\cpuregs[12] [8]), .B1 (n_484), .Y (n_4416));
  AOI22X1 g176697(.A0 (\cpuregs[20] [8]), .A1 (n_488), .B0
       (\cpuregs[23] [8]), .B1 (n_464), .Y (n_4415));
  AOI22X1 g176698(.A0 (\cpuregs[16] [8]), .A1 (n_478), .B0
       (\cpuregs[21] [8]), .B1 (n_468), .Y (n_4414));
  AOI22X1 g176699(.A0 (\cpuregs[17] [8]), .A1 (n_486), .B0
       (\cpuregs[18] [8]), .B1 (n_492), .Y (n_4413));
  AOI22X1 g176700(.A0 (\cpuregs[26] [8]), .A1 (n_490), .B0
       (\cpuregs[27] [8]), .B1 (n_498), .Y (n_4412));
  AOI22X1 g176701(.A0 (\cpuregs[28] [8]), .A1 (n_480), .B0
       (\cpuregs[29] [8]), .B1 (n_458), .Y (n_4411));
  AOI22X1 g176702(.A0 (\cpuregs[30] [8]), .A1 (n_500), .B0
       (\cpuregs[31] [8]), .B1 (n_476), .Y (n_4410));
  AOI22X1 g176703(.A0 (\cpuregs[24] [8]), .A1 (n_494), .B0
       (\cpuregs[25] [8]), .B1 (n_496), .Y (n_4409));
  AOI22X1 g176704(.A0 (\cpuregs[3] [9]), .A1 (n_423), .B0
       (\cpuregs[15] [9]), .B1 (n_462), .Y (n_4408));
  AOI22X1 g176705(.A0 (\cpuregs[1] [9]), .A1 (n_456), .B0
       (\cpuregs[2] [9]), .B1 (n_425), .Y (n_4407));
  AOI22X1 g176706(.A0 (\cpuregs[4] [9]), .A1 (n_424), .B0
       (\cpuregs[6] [9]), .B1 (n_333), .Y (n_4406));
  AOI22X1 g176707(.A0 (\cpuregs[13] [9]), .A1 (n_454), .B0
       (\cpuregs[14] [9]), .B1 (n_450), .Y (n_4405));
  AOI22X1 g176708(.A0 (\cpuregs[8] [9]), .A1 (n_466), .B0
       (\cpuregs[7] [9]), .B1 (n_474), .Y (n_4404));
  AOI22X1 g176709(.A0 (\cpuregs[10] [9]), .A1 (n_452), .B0
       (\cpuregs[11] [9]), .B1 (n_448), .Y (n_4403));
  AOI22X1 g176710(.A0 (\cpuregs[9] [9]), .A1 (n_470), .B0
       (\cpuregs[12] [9]), .B1 (n_484), .Y (n_4402));
  AOI22X1 g176711(.A0 (\cpuregs[16] [9]), .A1 (n_478), .B0
       (\cpuregs[23] [9]), .B1 (n_464), .Y (n_4401));
  AOI22X1 g176712(.A0 (\cpuregs[17] [9]), .A1 (n_486), .B0
       (\cpuregs[18] [9]), .B1 (n_492), .Y (n_4400));
  AOI22X1 g176713(.A0 (\cpuregs[20] [9]), .A1 (n_488), .B0
       (\cpuregs[19] [9]), .B1 (n_502), .Y (n_4399));
  AOI22X1 g176714(.A0 (\cpuregs[30] [9]), .A1 (n_500), .B0
       (\cpuregs[31] [9]), .B1 (n_476), .Y (n_4398));
  AOI22X1 g176715(.A0 (\cpuregs[28] [9]), .A1 (n_480), .B0
       (\cpuregs[29] [9]), .B1 (n_458), .Y (n_4397));
  AOI22X1 g176716(.A0 (\cpuregs[26] [9]), .A1 (n_490), .B0
       (\cpuregs[27] [9]), .B1 (n_498), .Y (n_4396));
  AOI22X1 g176717(.A0 (\cpuregs[24] [9]), .A1 (n_494), .B0
       (\cpuregs[25] [9]), .B1 (n_496), .Y (n_4395));
  AOI22X1 g176718(.A0 (\cpuregs[9] [10]), .A1 (n_470), .B0
       (\cpuregs[10] [10]), .B1 (n_452), .Y (n_4394));
  AOI22X1 g176719(.A0 (\cpuregs[8] [10]), .A1 (n_466), .B0
       (\cpuregs[7] [10]), .B1 (n_474), .Y (n_4393));
  AO22X1 g176720(.A0 (\cpuregs[11] [10]), .A1 (n_448), .B0
       (\cpuregs[14] [10]), .B1 (n_450), .Y (n_4392));
  AOI22X1 g176721(.A0 (\cpuregs[5] [10]), .A1 (n_291), .B0
       (\cpuregs[3] [10]), .B1 (n_423), .Y (n_4391));
  AOI22X1 g176722(.A0 (\cpuregs[26] [10]), .A1 (n_490), .B0
       (\cpuregs[29] [10]), .B1 (n_458), .Y (n_4390));
  AOI22X1 g176723(.A0 (\cpuregs[25] [10]), .A1 (n_496), .B0
       (\cpuregs[28] [10]), .B1 (n_480), .Y (n_4389));
  AOI22X1 g176724(.A0 (\cpuregs[27] [10]), .A1 (n_498), .B0
       (\cpuregs[30] [10]), .B1 (n_500), .Y (n_4388));
  AOI22X1 g176725(.A0 (\cpuregs[18] [10]), .A1 (n_492), .B0
       (\cpuregs[19] [10]), .B1 (n_502), .Y (n_4387));
  AOI22X1 g176726(.A0 (\cpuregs[20] [10]), .A1 (n_488), .B0
       (\cpuregs[21] [10]), .B1 (n_468), .Y (n_4386));
  AOI22X1 g176727(.A0 (\cpuregs[22] [10]), .A1 (n_482), .B0
       (\cpuregs[23] [10]), .B1 (n_464), .Y (n_4385));
  AOI22X1 g176728(.A0 (\cpuregs[16] [10]), .A1 (n_478), .B0
       (\cpuregs[17] [10]), .B1 (n_486), .Y (n_4384));
  AOI22X1 g176729(.A0 (\cpuregs[3] [11]), .A1 (n_423), .B0
       (\cpuregs[15] [11]), .B1 (n_462), .Y (n_4383));
  AOI22X1 g176730(.A0 (\cpuregs[1] [11]), .A1 (n_456), .B0
       (\cpuregs[2] [11]), .B1 (n_425), .Y (n_4382));
  AOI22X1 g176731(.A0 (\cpuregs[4] [11]), .A1 (n_424), .B0
       (\cpuregs[6] [11]), .B1 (n_333), .Y (n_4381));
  AOI22X1 g176732(.A0 (\cpuregs[13] [11]), .A1 (n_454), .B0
       (\cpuregs[14] [11]), .B1 (n_450), .Y (n_4380));
  AOI22X1 g176733(.A0 (\cpuregs[8] [11]), .A1 (n_466), .B0
       (\cpuregs[7] [11]), .B1 (n_474), .Y (n_4379));
  AOI22X1 g176734(.A0 (\cpuregs[10] [11]), .A1 (n_452), .B0
       (\cpuregs[11] [11]), .B1 (n_448), .Y (n_4378));
  AOI22X1 g176735(.A0 (\cpuregs[9] [11]), .A1 (n_470), .B0
       (\cpuregs[12] [11]), .B1 (n_484), .Y (n_4377));
  AOI22X1 g176736(.A0 (\cpuregs[20] [11]), .A1 (n_488), .B0
       (\cpuregs[19] [11]), .B1 (n_502), .Y (n_4376));
  AOI22X1 g176737(.A0 (\cpuregs[16] [11]), .A1 (n_478), .B0
       (\cpuregs[21] [11]), .B1 (n_468), .Y (n_4375));
  AOI22X1 g176738(.A0 (\cpuregs[17] [11]), .A1 (n_486), .B0
       (\cpuregs[22] [11]), .B1 (n_482), .Y (n_4374));
  AOI22X1 g176739(.A0 (\cpuregs[30] [11]), .A1 (n_500), .B0
       (\cpuregs[31] [11]), .B1 (n_476), .Y (n_4373));
  AOI22X1 g176740(.A0 (\cpuregs[26] [11]), .A1 (n_490), .B0
       (\cpuregs[27] [11]), .B1 (n_498), .Y (n_4372));
  AOI22X1 g176741(.A0 (\cpuregs[28] [11]), .A1 (n_480), .B0
       (\cpuregs[29] [11]), .B1 (n_458), .Y (n_4371));
  AOI22X1 g176742(.A0 (\cpuregs[24] [11]), .A1 (n_494), .B0
       (\cpuregs[25] [11]), .B1 (n_496), .Y (n_4370));
  AOI22X1 g176743(.A0 (\cpuregs[3] [12]), .A1 (n_423), .B0
       (\cpuregs[15] [12]), .B1 (n_462), .Y (n_4369));
  AOI22X1 g176744(.A0 (\cpuregs[1] [12]), .A1 (n_456), .B0
       (\cpuregs[2] [12]), .B1 (n_425), .Y (n_4368));
  AOI22X1 g176745(.A0 (\cpuregs[4] [12]), .A1 (n_424), .B0
       (\cpuregs[6] [12]), .B1 (n_333), .Y (n_4367));
  AOI22X1 g176746(.A0 (\cpuregs[9] [12]), .A1 (n_470), .B0
       (\cpuregs[13] [12]), .B1 (n_454), .Y (n_4366));
  AOI22X1 g176747(.A0 (\cpuregs[10] [12]), .A1 (n_452), .B0
       (\cpuregs[14] [12]), .B1 (n_450), .Y (n_4365));
  AOI22X1 g176748(.A0 (\cpuregs[12] [12]), .A1 (n_484), .B0
       (\cpuregs[11] [12]), .B1 (n_448), .Y (n_4364));
  AOI22X1 g176749(.A0 (\cpuregs[8] [12]), .A1 (n_466), .B0
       (\cpuregs[7] [12]), .B1 (n_474), .Y (n_4363));
  AOI22X1 g176750(.A0 (\cpuregs[25] [12]), .A1 (n_496), .B0
       (\cpuregs[30] [12]), .B1 (n_500), .Y (n_4362));
  AOI22X1 g176751(.A0 (\cpuregs[24] [12]), .A1 (n_494), .B0
       (\cpuregs[27] [12]), .B1 (n_498), .Y (n_4361));
  AOI22X1 g176752(.A0 (\cpuregs[28] [12]), .A1 (n_480), .B0
       (\cpuregs[31] [12]), .B1 (n_476), .Y (n_4360));
  AOI22X1 g176753(.A0 (\cpuregs[18] [12]), .A1 (n_492), .B0
       (\cpuregs[19] [12]), .B1 (n_502), .Y (n_4359));
  AOI22X1 g176754(.A0 (\cpuregs[20] [12]), .A1 (n_488), .B0
       (\cpuregs[21] [12]), .B1 (n_468), .Y (n_4358));
  AOI22X1 g176755(.A0 (\cpuregs[22] [12]), .A1 (n_482), .B0
       (\cpuregs[23] [12]), .B1 (n_464), .Y (n_4357));
  AOI22X1 g176756(.A0 (\cpuregs[16] [12]), .A1 (n_478), .B0
       (\cpuregs[17] [12]), .B1 (n_486), .Y (n_4356));
  AOI22X1 g176757(.A0 (\cpuregs[13] [13]), .A1 (n_454), .B0
       (\cpuregs[14] [13]), .B1 (n_450), .Y (n_4355));
  AOI22X1 g176758(.A0 (\cpuregs[9] [13]), .A1 (n_470), .B0
       (\cpuregs[10] [13]), .B1 (n_452), .Y (n_4354));
  AO22X1 g176759(.A0 (\cpuregs[8] [13]), .A1 (n_466), .B0
       (\cpuregs[12] [13]), .B1 (n_484), .Y (n_4353));
  AOI22X1 g176760(.A0 (\cpuregs[3] [13]), .A1 (n_423), .B0
       (\cpuregs[6] [13]), .B1 (n_333), .Y (n_4352));
  AOI22X1 g176761(.A0 (\cpuregs[26] [13]), .A1 (n_490), .B0
       (\cpuregs[29] [13]), .B1 (n_458), .Y (n_4351));
  AOI22X1 g176762(.A0 (\cpuregs[25] [13]), .A1 (n_496), .B0
       (\cpuregs[28] [13]), .B1 (n_480), .Y (n_4350));
  AOI22X1 g176763(.A0 (\cpuregs[27] [13]), .A1 (n_498), .B0
       (\cpuregs[30] [13]), .B1 (n_500), .Y (n_4349));
  AOI22X1 g176764(.A0 (\cpuregs[22] [13]), .A1 (n_482), .B0
       (\cpuregs[23] [13]), .B1 (n_464), .Y (n_4348));
  AOI22X1 g176765(.A0 (\cpuregs[20] [13]), .A1 (n_488), .B0
       (\cpuregs[21] [13]), .B1 (n_468), .Y (n_4347));
  AOI22X1 g176766(.A0 (\cpuregs[18] [13]), .A1 (n_492), .B0
       (\cpuregs[19] [13]), .B1 (n_502), .Y (n_4346));
  AOI22X1 g176767(.A0 (\cpuregs[16] [13]), .A1 (n_478), .B0
       (\cpuregs[17] [13]), .B1 (n_486), .Y (n_4345));
  AO22X1 g176768(.A0 (\cpuregs[4] [14]), .A1 (n_424), .B0
       (\cpuregs[5] [14]), .B1 (n_291), .Y (n_4344));
  AOI22X1 g176769(.A0 (\cpuregs[15] [14]), .A1 (n_462), .B0 (n_833),
       .B1 (n_66), .Y (n_4343));
  AOI22X1 g176770(.A0 (\cpuregs[1] [14]), .A1 (n_456), .B0
       (reg_pc[14]), .B1 (n_961), .Y (n_4342));
  AOI22X1 g176771(.A0 (\cpuregs[7] [14]), .A1 (n_474), .B0
       (\cpuregs[14] [14]), .B1 (n_450), .Y (n_4341));
  AOI22X1 g176772(.A0 (\cpuregs[8] [14]), .A1 (n_466), .B0
       (\cpuregs[13] [14]), .B1 (n_454), .Y (n_4340));
  AOI22X1 g176773(.A0 (\cpuregs[12] [14]), .A1 (n_484), .B0
       (\cpuregs[11] [14]), .B1 (n_448), .Y (n_4339));
  AOI22X1 g176774(.A0 (\cpuregs[9] [14]), .A1 (n_470), .B0
       (\cpuregs[10] [14]), .B1 (n_452), .Y (n_4338));
  AOI22X1 g176775(.A0 (\cpuregs[30] [14]), .A1 (n_500), .B0
       (\cpuregs[31] [14]), .B1 (n_476), .Y (n_4337));
  AOI22X1 g176776(.A0 (\cpuregs[26] [14]), .A1 (n_490), .B0
       (\cpuregs[27] [14]), .B1 (n_498), .Y (n_4336));
  AOI22X1 g176777(.A0 (\cpuregs[28] [14]), .A1 (n_480), .B0
       (\cpuregs[29] [14]), .B1 (n_458), .Y (n_4335));
  AOI22X1 g176778(.A0 (\cpuregs[24] [14]), .A1 (n_494), .B0
       (\cpuregs[25] [14]), .B1 (n_496), .Y (n_4334));
  AOI22X1 g176779(.A0 (\cpuregs[18] [14]), .A1 (n_492), .B0
       (\cpuregs[19] [14]), .B1 (n_502), .Y (n_4333));
  AOI22X1 g176780(.A0 (\cpuregs[20] [14]), .A1 (n_488), .B0
       (\cpuregs[21] [14]), .B1 (n_468), .Y (n_4332));
  AOI22X1 g176781(.A0 (\cpuregs[22] [14]), .A1 (n_482), .B0
       (\cpuregs[23] [14]), .B1 (n_464), .Y (n_4331));
  AOI22X1 g176782(.A0 (\cpuregs[16] [14]), .A1 (n_478), .B0
       (\cpuregs[17] [14]), .B1 (n_486), .Y (n_4330));
  AOI22X1 g176783(.A0 (\cpuregs[20] [15]), .A1 (n_488), .B0
       (\cpuregs[21] [15]), .B1 (n_468), .Y (n_4329));
  AOI22X1 g176784(.A0 (\cpuregs[16] [15]), .A1 (n_478), .B0
       (\cpuregs[17] [15]), .B1 (n_486), .Y (n_4328));
  AO22X1 g176785(.A0 (\cpuregs[22] [15]), .A1 (n_482), .B0
       (\cpuregs[23] [15]), .B1 (n_464), .Y (n_4327));
  AOI22X1 g176786(.A0 (\cpuregs[26] [15]), .A1 (n_490), .B0
       (\cpuregs[27] [15]), .B1 (n_498), .Y (n_4326));
  AOI22X1 g176787(.A0 (\cpuregs[28] [15]), .A1 (n_480), .B0
       (\cpuregs[29] [15]), .B1 (n_458), .Y (n_4325));
  AOI22X1 g176788(.A0 (\cpuregs[30] [15]), .A1 (n_500), .B0
       (\cpuregs[31] [15]), .B1 (n_476), .Y (n_4324));
  AOI22X1 g176789(.A0 (\cpuregs[24] [15]), .A1 (n_494), .B0
       (\cpuregs[25] [15]), .B1 (n_496), .Y (n_4323));
  AOI22X1 g176790(.A0 (\cpuregs[4] [15]), .A1 (n_424), .B0
       (\cpuregs[3] [15]), .B1 (n_423), .Y (n_4322));
  AOI22X1 g176791(.A0 (\cpuregs[5] [15]), .A1 (n_291), .B0
       (\cpuregs[6] [15]), .B1 (n_333), .Y (n_4321));
  AOI22X1 g176792(.A0 (\cpuregs[7] [15]), .A1 (n_474), .B0
       (\cpuregs[14] [15]), .B1 (n_450), .Y (n_4320));
  AOI22X1 g176793(.A0 (\cpuregs[8] [15]), .A1 (n_466), .B0
       (\cpuregs[13] [15]), .B1 (n_454), .Y (n_4319));
  AOI22X1 g176794(.A0 (\cpuregs[12] [15]), .A1 (n_484), .B0
       (\cpuregs[11] [15]), .B1 (n_448), .Y (n_4318));
  AOI22X1 g176795(.A0 (\cpuregs[9] [15]), .A1 (n_470), .B0
       (\cpuregs[10] [15]), .B1 (n_452), .Y (n_4317));
  AOI22X1 g176796(.A0 (\cpuregs[5] [16]), .A1 (n_291), .B0
       (\cpuregs[15] [16]), .B1 (n_462), .Y (n_4316));
  AOI22X1 g176797(.A0 (\cpuregs[4] [16]), .A1 (n_424), .B0
       (\cpuregs[6] [16]), .B1 (n_333), .Y (n_4315));
  AOI22X1 g176798(.A0 (\cpuregs[13] [16]), .A1 (n_454), .B0
       (\cpuregs[14] [16]), .B1 (n_450), .Y (n_4314));
  AOI22X1 g176799(.A0 (\cpuregs[12] [16]), .A1 (n_484), .B0
       (\cpuregs[11] [16]), .B1 (n_448), .Y (n_4313));
  AOI22X1 g176800(.A0 (\cpuregs[10] [16]), .A1 (n_452), .B0
       (\cpuregs[7] [16]), .B1 (n_474), .Y (n_4312));
  AOI22X1 g176801(.A0 (\cpuregs[8] [16]), .A1 (n_466), .B0
       (\cpuregs[9] [16]), .B1 (n_470), .Y (n_4311));
  AOI22X1 g176802(.A0 (\cpuregs[30] [16]), .A1 (n_500), .B0
       (\cpuregs[31] [16]), .B1 (n_476), .Y (n_4310));
  AOI22X1 g176803(.A0 (\cpuregs[26] [16]), .A1 (n_490), .B0
       (\cpuregs[27] [16]), .B1 (n_498), .Y (n_4309));
  AOI22X1 g176804(.A0 (\cpuregs[28] [16]), .A1 (n_480), .B0
       (\cpuregs[29] [16]), .B1 (n_458), .Y (n_4308));
  AOI22X1 g176805(.A0 (\cpuregs[24] [16]), .A1 (n_494), .B0
       (\cpuregs[25] [16]), .B1 (n_496), .Y (n_4307));
  AOI22X1 g176806(.A0 (\cpuregs[18] [16]), .A1 (n_492), .B0
       (\cpuregs[19] [16]), .B1 (n_502), .Y (n_4306));
  AOI22X1 g176807(.A0 (\cpuregs[20] [16]), .A1 (n_488), .B0
       (\cpuregs[21] [16]), .B1 (n_468), .Y (n_4305));
  AOI22X1 g176808(.A0 (\cpuregs[22] [16]), .A1 (n_482), .B0
       (\cpuregs[23] [16]), .B1 (n_464), .Y (n_4304));
  AOI22X1 g176809(.A0 (\cpuregs[16] [16]), .A1 (n_478), .B0
       (\cpuregs[17] [16]), .B1 (n_486), .Y (n_4303));
  AOI22X1 g176810(.A0 (\cpuregs[3] [17]), .A1 (n_423), .B0
       (\cpuregs[15] [17]), .B1 (n_462), .Y (n_4302));
  AOI22X1 g176811(.A0 (\cpuregs[1] [17]), .A1 (n_456), .B0
       (\cpuregs[2] [17]), .B1 (n_425), .Y (n_4301));
  AOI22X1 g176812(.A0 (\cpuregs[4] [17]), .A1 (n_424), .B0
       (\cpuregs[6] [17]), .B1 (n_333), .Y (n_4300));
  AOI22X1 g176813(.A0 (\cpuregs[8] [17]), .A1 (n_466), .B0
       (\cpuregs[7] [17]), .B1 (n_474), .Y (n_4299));
  AOI22X1 g176814(.A0 (\cpuregs[13] [17]), .A1 (n_454), .B0
       (\cpuregs[14] [17]), .B1 (n_450), .Y (n_4298));
  AOI22X1 g176815(.A0 (\cpuregs[10] [17]), .A1 (n_452), .B0
       (\cpuregs[11] [17]), .B1 (n_448), .Y (n_4297));
  AOI22X1 g176816(.A0 (\cpuregs[9] [17]), .A1 (n_470), .B0
       (\cpuregs[12] [17]), .B1 (n_484), .Y (n_4296));
  AOI22X1 g176817(.A0 (\cpuregs[28] [17]), .A1 (n_480), .B0
       (\cpuregs[27] [17]), .B1 (n_498), .Y (n_4295));
  AOI22X1 g176818(.A0 (\cpuregs[24] [17]), .A1 (n_494), .B0
       (\cpuregs[29] [17]), .B1 (n_458), .Y (n_4294));
  AOI22X1 g176819(.A0 (\cpuregs[25] [17]), .A1 (n_496), .B0
       (\cpuregs[30] [17]), .B1 (n_500), .Y (n_4293));
  AOI22X1 g176820(.A0 (\cpuregs[22] [17]), .A1 (n_482), .B0
       (\cpuregs[23] [17]), .B1 (n_464), .Y (n_4292));
  AOI22X1 g176821(.A0 (\cpuregs[20] [17]), .A1 (n_488), .B0
       (\cpuregs[21] [17]), .B1 (n_468), .Y (n_4291));
  OAI21X1 g176822(.A0 (n_2440), .A1 (n_1), .B0 (n_1330), .Y (n_4712));
  NOR4BBX1 g176993(.AN (n_3250), .BN (n_2511), .C (n_3043), .D
       (n_3466), .Y (n_296));
  INVX1 g176999(.A (n_4289), .Y (n_4290));
  MX2X1 g177000(.A (n_376), .B (\cpuregs[13] [25]), .S0 (n_3233), .Y
       (n_4282));
  MX2X1 g177001(.A (n_396), .B (\cpuregs[5] [16]), .S0 (n_3221), .Y
       (n_4281));
  MX2X1 g177002(.A (n_414), .B (\cpuregs[5] [15]), .S0 (n_3221), .Y
       (n_4280));
  MX2X1 g177003(.A (n_374), .B (\cpuregs[5] [14]), .S0 (n_3221), .Y
       (n_4279));
  MX2X1 g177004(.A (n_388), .B (\cpuregs[5] [13]), .S0 (n_3221), .Y
       (n_4278));
  MX2X1 g177005(.A (n_384), .B (\cpuregs[5] [12]), .S0 (n_3221), .Y
       (n_4277));
  MX2X1 g177006(.A (n_402), .B (\cpuregs[5] [11]), .S0 (n_3221), .Y
       (n_4276));
  MX2X1 g177007(.A (n_408), .B (\cpuregs[5] [10]), .S0 (n_3221), .Y
       (n_4275));
  MX2X1 g177008(.A (n_372), .B (\cpuregs[5] [9]), .S0 (n_3221), .Y
       (n_4274));
  MX2X1 g177009(.A (n_418), .B (\cpuregs[5] [8]), .S0 (n_3221), .Y
       (n_4273));
  MX2X1 g177010(.A (n_386), .B (\cpuregs[5] [7]), .S0 (n_3221), .Y
       (n_4272));
  MX2X1 g177011(.A (n_362), .B (\cpuregs[5] [6]), .S0 (n_3221), .Y
       (n_4271));
  MX2X1 g177012(.A (n_394), .B (\cpuregs[5] [5]), .S0 (n_3221), .Y
       (n_4270));
  MX2X1 g177013(.A (n_416), .B (\cpuregs[5] [4]), .S0 (n_3221), .Y
       (n_4269));
  MX2X1 g177014(.A (n_368), .B (\cpuregs[5] [3]), .S0 (n_3221), .Y
       (n_4268));
  MX2X1 g177015(.A (n_366), .B (\cpuregs[5] [2]), .S0 (n_3221), .Y
       (n_4267));
  MX2X1 g177016(.A (n_398), .B (\cpuregs[5] [1]), .S0 (n_3221), .Y
       (n_4266));
  MX2X1 g177017(.A (n_398), .B (\cpuregs[6] [1]), .S0 (n_3215), .Y
       (n_4265));
  MX2X1 g177018(.A (n_366), .B (\cpuregs[6] [2]), .S0 (n_3215), .Y
       (n_4264));
  MX2X1 g177019(.A (n_404), .B (\cpuregs[22] [31]), .S0 (n_3213), .Y
       (n_4263));
  MX2X1 g177020(.A (n_370), .B (\cpuregs[22] [30]), .S0 (n_3213), .Y
       (n_4262));
  MX2X1 g177021(.A (n_392), .B (\cpuregs[22] [29]), .S0 (n_3213), .Y
       (n_4261));
  MX2X1 g177022(.A (n_390), .B (\cpuregs[22] [28]), .S0 (n_3213), .Y
       (n_4260));
  MX2X1 g177023(.A (n_406), .B (\cpuregs[22] [27]), .S0 (n_3213), .Y
       (n_4259));
  MX2X1 g177024(.A (n_400), .B (\cpuregs[22] [26]), .S0 (n_3213), .Y
       (n_4258));
  MX2X1 g177025(.A (n_376), .B (\cpuregs[22] [25]), .S0 (n_3213), .Y
       (n_4257));
  MX2X1 g177026(.A (n_378), .B (\cpuregs[22] [24]), .S0 (n_3213), .Y
       (n_4256));
  MX2X1 g177027(.A (n_380), .B (\cpuregs[22] [23]), .S0 (n_3213), .Y
       (n_4255));
  MX2X1 g177028(.A (n_1513), .B (\cpuregs[22] [22]), .S0 (n_3213), .Y
       (n_4254));
  MX2X1 g177029(.A (n_1515), .B (\cpuregs[22] [21]), .S0 (n_3213), .Y
       (n_4253));
  MX2X1 g177030(.A (n_364), .B (\cpuregs[22] [20]), .S0 (n_3213), .Y
       (n_4252));
  MX2X1 g177031(.A (n_1518), .B (\cpuregs[22] [19]), .S0 (n_3213), .Y
       (n_4251));
  MX2X1 g177032(.A (n_382), .B (\cpuregs[22] [18]), .S0 (n_3213), .Y
       (n_4250));
  MX2X1 g177033(.A (n_412), .B (\cpuregs[22] [17]), .S0 (n_3213), .Y
       (n_4249));
  MX2X1 g177034(.A (n_396), .B (\cpuregs[22] [16]), .S0 (n_3213), .Y
       (n_4248));
  MX2X1 g177035(.A (n_414), .B (\cpuregs[22] [15]), .S0 (n_3213), .Y
       (n_4247));
  MX2X1 g177036(.A (n_374), .B (\cpuregs[22] [14]), .S0 (n_3213), .Y
       (n_4246));
  MX2X1 g177037(.A (n_388), .B (\cpuregs[22] [13]), .S0 (n_3213), .Y
       (n_4245));
  MX2X1 g177038(.A (n_384), .B (\cpuregs[22] [12]), .S0 (n_3213), .Y
       (n_4244));
  MX2X1 g177039(.A (n_402), .B (\cpuregs[22] [11]), .S0 (n_3213), .Y
       (n_4243));
  MX2X1 g177040(.A (n_408), .B (\cpuregs[22] [10]), .S0 (n_3213), .Y
       (n_4242));
  MX2X1 g177041(.A (n_372), .B (\cpuregs[22] [9]), .S0 (n_3213), .Y
       (n_4241));
  MX2X1 g177042(.A (n_418), .B (\cpuregs[22] [8]), .S0 (n_3213), .Y
       (n_4240));
  MX2X1 g177043(.A (n_386), .B (\cpuregs[22] [7]), .S0 (n_3213), .Y
       (n_4239));
  MX2X1 g177044(.A (n_362), .B (\cpuregs[22] [6]), .S0 (n_3213), .Y
       (n_4238));
  MX2X1 g177045(.A (n_394), .B (\cpuregs[22] [5]), .S0 (n_3213), .Y
       (n_4237));
  MX2X1 g177046(.A (n_416), .B (\cpuregs[22] [4]), .S0 (n_3213), .Y
       (n_4236));
  MX2X1 g177047(.A (n_368), .B (\cpuregs[22] [3]), .S0 (n_3213), .Y
       (n_4235));
  MX2X1 g177048(.A (n_366), .B (\cpuregs[22] [2]), .S0 (n_3213), .Y
       (n_4234));
  MX2X1 g177049(.A (n_398), .B (\cpuregs[22] [1]), .S0 (n_3213), .Y
       (n_4233));
  MX2X1 g177050(.A (n_404), .B (\cpuregs[3] [31]), .S0 (n_3219), .Y
       (n_4232));
  MX2X1 g177051(.A (n_404), .B (\cpuregs[21] [31]), .S0 (n_3214), .Y
       (n_4231));
  MX2X1 g177052(.A (n_370), .B (\cpuregs[3] [30]), .S0 (n_3219), .Y
       (n_4230));
  MX2X1 g177053(.A (n_370), .B (\cpuregs[21] [30]), .S0 (n_3214), .Y
       (n_4229));
  MX2X1 g177054(.A (n_392), .B (\cpuregs[21] [29]), .S0 (n_3214), .Y
       (n_4228));
  MX2X1 g177055(.A (n_392), .B (\cpuregs[3] [29]), .S0 (n_3219), .Y
       (n_4227));
  MX2X1 g177056(.A (n_390), .B (\cpuregs[3] [28]), .S0 (n_3219), .Y
       (n_4226));
  MX2X1 g177057(.A (n_390), .B (\cpuregs[21] [28]), .S0 (n_3214), .Y
       (n_4225));
  MX2X1 g177058(.A (n_406), .B (\cpuregs[21] [27]), .S0 (n_3214), .Y
       (n_4224));
  MX2X1 g177059(.A (n_400), .B (\cpuregs[21] [26]), .S0 (n_3214), .Y
       (n_4223));
  MX2X1 g177060(.A (n_406), .B (\cpuregs[3] [27]), .S0 (n_3219), .Y
       (n_4222));
  MX2X1 g177061(.A (n_376), .B (\cpuregs[21] [25]), .S0 (n_3214), .Y
       (n_4221));
  MX2X1 g177062(.A (n_378), .B (\cpuregs[21] [24]), .S0 (n_3214), .Y
       (n_4220));
  MX2X1 g177063(.A (n_380), .B (\cpuregs[21] [23]), .S0 (n_3214), .Y
       (n_4219));
  MX2X1 g177064(.A (n_400), .B (\cpuregs[3] [26]), .S0 (n_3219), .Y
       (n_4218));
  MX2X1 g177065(.A (n_378), .B (\cpuregs[3] [24]), .S0 (n_3219), .Y
       (n_4217));
  MX2X1 g177066(.A (n_1513), .B (\cpuregs[21] [22]), .S0 (n_3214), .Y
       (n_4216));
  MX2X1 g177067(.A (n_1515), .B (\cpuregs[21] [21]), .S0 (n_3214), .Y
       (n_4215));
  MX2X1 g177068(.A (n_376), .B (\cpuregs[3] [25]), .S0 (n_3219), .Y
       (n_4214));
  MX2X1 g177069(.A (n_364), .B (\cpuregs[21] [20]), .S0 (n_3214), .Y
       (n_4213));
  MX2X1 g177070(.A (n_1518), .B (\cpuregs[21] [19]), .S0 (n_3214), .Y
       (n_4212));
  MX2X1 g177071(.A (n_382), .B (\cpuregs[21] [18]), .S0 (n_3214), .Y
       (n_4211));
  MX2X1 g177072(.A (n_412), .B (\cpuregs[21] [17]), .S0 (n_3214), .Y
       (n_4210));
  MX2X1 g177073(.A (n_380), .B (\cpuregs[3] [23]), .S0 (n_3219), .Y
       (n_4209));
  MX2X1 g177074(.A (n_396), .B (\cpuregs[21] [16]), .S0 (n_3214), .Y
       (n_4208));
  MX2X1 g177075(.A (n_414), .B (\cpuregs[21] [15]), .S0 (n_3214), .Y
       (n_4207));
  OAI22X1 g177076(.A0 (n_3219), .A1 (n_1512), .B0 (n_606), .B1 (n_697),
       .Y (n_4206));
  MX2X1 g177077(.A (n_374), .B (\cpuregs[21] [14]), .S0 (n_3214), .Y
       (n_4205));
  MX2X1 g177078(.A (n_388), .B (\cpuregs[21] [13]), .S0 (n_3214), .Y
       (n_4204));
  OAI22X1 g177079(.A0 (n_3219), .A1 (n_1514), .B0 (n_655), .B1 (n_697),
       .Y (n_4203));
  MX2X1 g177080(.A (n_384), .B (\cpuregs[21] [12]), .S0 (n_3214), .Y
       (n_4202));
  MX2X1 g177081(.A (n_402), .B (\cpuregs[21] [11]), .S0 (n_3214), .Y
       (n_4201));
  MX2X1 g177082(.A (n_364), .B (\cpuregs[3] [20]), .S0 (n_3219), .Y
       (n_4200));
  MX2X1 g177083(.A (n_408), .B (\cpuregs[21] [10]), .S0 (n_3214), .Y
       (n_4199));
  MX2X1 g177084(.A (n_372), .B (\cpuregs[21] [9]), .S0 (n_3214), .Y
       (n_4198));
  MX2X1 g177085(.A (n_418), .B (\cpuregs[21] [8]), .S0 (n_3214), .Y
       (n_4197));
  OAI22X1 g177086(.A0 (n_3219), .A1 (n_1517), .B0 (n_604), .B1 (n_697),
       .Y (n_4196));
  MX2X1 g177087(.A (n_386), .B (\cpuregs[21] [7]), .S0 (n_3214), .Y
       (n_4195));
  MX2X1 g177088(.A (n_382), .B (\cpuregs[3] [18]), .S0 (n_3219), .Y
       (n_4194));
  MX2X1 g177089(.A (n_362), .B (\cpuregs[21] [6]), .S0 (n_3214), .Y
       (n_4193));
  MX2X1 g177090(.A (n_412), .B (\cpuregs[3] [17]), .S0 (n_3219), .Y
       (n_4192));
  MX2X1 g177091(.A (n_398), .B (\cpuregs[27] [1]), .S0 (n_3220), .Y
       (n_4191));
  MX2X1 g177092(.A (n_394), .B (\cpuregs[21] [5]), .S0 (n_3214), .Y
       (n_4190));
  MX2X1 g177093(.A (n_416), .B (\cpuregs[21] [4]), .S0 (n_3214), .Y
       (n_4189));
  MX2X1 g177094(.A (n_396), .B (\cpuregs[3] [16]), .S0 (n_3219), .Y
       (n_4188));
  MX2X1 g177095(.A (n_368), .B (\cpuregs[21] [3]), .S0 (n_3214), .Y
       (n_4187));
  MX2X1 g177096(.A (n_366), .B (\cpuregs[21] [2]), .S0 (n_3214), .Y
       (n_4186));
  MX2X1 g177097(.A (n_398), .B (\cpuregs[21] [1]), .S0 (n_3214), .Y
       (n_4185));
  MX2X1 g177098(.A (n_414), .B (\cpuregs[3] [15]), .S0 (n_3219), .Y
       (n_4184));
  MX2X1 g177099(.A (n_374), .B (\cpuregs[3] [14]), .S0 (n_3219), .Y
       (n_4183));
  MX2X1 g177100(.A (n_368), .B (\cpuregs[27] [3]), .S0 (n_3220), .Y
       (n_4182));
  MX2X1 g177101(.A (n_388), .B (\cpuregs[3] [13]), .S0 (n_3219), .Y
       (n_4181));
  MX2X1 g177102(.A (n_384), .B (\cpuregs[3] [12]), .S0 (n_3219), .Y
       (n_4180));
  MX2X1 g177103(.A (n_402), .B (\cpuregs[3] [11]), .S0 (n_3219), .Y
       (n_4179));
  MX2X1 g177104(.A (n_408), .B (\cpuregs[3] [10]), .S0 (n_3219), .Y
       (n_4178));
  MX2X1 g177105(.A (n_372), .B (\cpuregs[3] [9]), .S0 (n_3219), .Y
       (n_4177));
  MX2X1 g177106(.A (n_418), .B (\cpuregs[3] [8]), .S0 (n_3219), .Y
       (n_4176));
  MX2X1 g177107(.A (n_416), .B (\cpuregs[3] [4]), .S0 (n_3219), .Y
       (n_4175));
  MX2X1 g177108(.A (n_386), .B (\cpuregs[3] [7]), .S0 (n_3219), .Y
       (n_4174));
  MX2X1 g177109(.A (n_372), .B (\cpuregs[27] [9]), .S0 (n_3220), .Y
       (n_4173));
  MX2X1 g177110(.A (n_362), .B (\cpuregs[3] [6]), .S0 (n_3219), .Y
       (n_4172));
  MX2X1 g177111(.A (n_394), .B (\cpuregs[3] [5]), .S0 (n_3219), .Y
       (n_4171));
  MX2X1 g177112(.A (n_368), .B (\cpuregs[3] [3]), .S0 (n_3219), .Y
       (n_4170));
  MX2X1 g177113(.A (n_366), .B (\cpuregs[3] [2]), .S0 (n_3219), .Y
       (n_4169));
  MX2X1 g177114(.A (n_398), .B (\cpuregs[3] [1]), .S0 (n_3219), .Y
       (n_4168));
  MX2X1 g177115(.A (n_404), .B (\cpuregs[19] [31]), .S0 (n_3216), .Y
       (n_4167));
  MX2X1 g177116(.A (n_404), .B (\cpuregs[2] [31]), .S0 (n_3218), .Y
       (n_4166));
  MX2X1 g177117(.A (n_370), .B (\cpuregs[19] [30]), .S0 (n_3216), .Y
       (n_4165));
  MX2X1 g177118(.A (n_370), .B (\cpuregs[2] [30]), .S0 (n_3218), .Y
       (n_4164));
  MX2X1 g177119(.A (n_392), .B (\cpuregs[19] [29]), .S0 (n_3216), .Y
       (n_4163));
  MX2X1 g177120(.A (n_390), .B (\cpuregs[19] [28]), .S0 (n_3216), .Y
       (n_4162));
  MX2X1 g177121(.A (n_392), .B (\cpuregs[2] [29]), .S0 (n_3218), .Y
       (n_4161));
  MX2X1 g177122(.A (n_406), .B (\cpuregs[19] [27]), .S0 (n_3216), .Y
       (n_4160));
  MX2X1 g177123(.A (n_400), .B (\cpuregs[19] [26]), .S0 (n_3216), .Y
       (n_4159));
  MX2X1 g177124(.A (n_376), .B (\cpuregs[19] [25]), .S0 (n_3216), .Y
       (n_4158));
  MX2X1 g177125(.A (n_390), .B (\cpuregs[2] [28]), .S0 (n_3218), .Y
       (n_4157));
  MX2X1 g177126(.A (n_378), .B (\cpuregs[19] [24]), .S0 (n_3216), .Y
       (n_4156));
  MX2X1 g177127(.A (n_406), .B (\cpuregs[2] [27]), .S0 (n_3218), .Y
       (n_4155));
  MX2X1 g177128(.A (n_380), .B (\cpuregs[19] [23]), .S0 (n_3216), .Y
       (n_4154));
  MX2X1 g177129(.A (n_378), .B (\cpuregs[2] [24]), .S0 (n_3218), .Y
       (n_4153));
  MX2X1 g177130(.A (n_1513), .B (\cpuregs[19] [22]), .S0 (n_3216), .Y
       (n_4152));
  MX2X1 g177131(.A (n_400), .B (\cpuregs[2] [26]), .S0 (n_3218), .Y
       (n_4151));
  MX2X1 g177132(.A (n_1515), .B (\cpuregs[19] [21]), .S0 (n_3216), .Y
       (n_4150));
  MX2X1 g177133(.A (n_364), .B (\cpuregs[19] [20]), .S0 (n_3216), .Y
       (n_4149));
  MX2X1 g177134(.A (n_1518), .B (\cpuregs[19] [19]), .S0 (n_3216), .Y
       (n_4148));
  MX2X1 g177135(.A (n_376), .B (\cpuregs[2] [25]), .S0 (n_3218), .Y
       (n_4147));
  MX2X1 g177136(.A (n_382), .B (\cpuregs[19] [18]), .S0 (n_3216), .Y
       (n_4146));
  MX2X1 g177137(.A (n_412), .B (\cpuregs[19] [17]), .S0 (n_3216), .Y
       (n_4145));
  MX2X1 g177138(.A (n_396), .B (\cpuregs[19] [16]), .S0 (n_3216), .Y
       (n_4144));
  MX2X1 g177139(.A (n_414), .B (\cpuregs[19] [15]), .S0 (n_3216), .Y
       (n_4143));
  MX2X1 g177140(.A (n_380), .B (\cpuregs[2] [23]), .S0 (n_3218), .Y
       (n_4142));
  MX2X1 g177141(.A (n_374), .B (\cpuregs[19] [14]), .S0 (n_3216), .Y
       (n_4141));
  MX2X1 g177142(.A (n_1513), .B (\cpuregs[2] [22]), .S0 (n_3218), .Y
       (n_4140));
  MX2X1 g177143(.A (n_1515), .B (\cpuregs[2] [21]), .S0 (n_3218), .Y
       (n_4139));
  MX2X1 g177144(.A (n_388), .B (\cpuregs[19] [13]), .S0 (n_3216), .Y
       (n_4138));
  MX2X1 g177145(.A (n_384), .B (\cpuregs[19] [12]), .S0 (n_3216), .Y
       (n_4137));
  MX2X1 g177146(.A (n_402), .B (\cpuregs[19] [11]), .S0 (n_3216), .Y
       (n_4136));
  MX2X1 g177147(.A (n_408), .B (\cpuregs[19] [10]), .S0 (n_3216), .Y
       (n_4135));
  MX2X1 g177148(.A (n_364), .B (\cpuregs[2] [20]), .S0 (n_3218), .Y
       (n_4134));
  MX2X1 g177149(.A (n_372), .B (\cpuregs[19] [9]), .S0 (n_3216), .Y
       (n_4133));
  MX2X1 g177150(.A (n_1518), .B (\cpuregs[2] [19]), .S0 (n_3218), .Y
       (n_4132));
  MX2X1 g177151(.A (n_418), .B (\cpuregs[19] [8]), .S0 (n_3216), .Y
       (n_4131));
  MX2X1 g177152(.A (n_382), .B (\cpuregs[2] [18]), .S0 (n_3218), .Y
       (n_4130));
  MX2X1 g177153(.A (n_386), .B (\cpuregs[19] [7]), .S0 (n_3216), .Y
       (n_4129));
  MX2X1 g177154(.A (n_362), .B (\cpuregs[19] [6]), .S0 (n_3216), .Y
       (n_4128));
  MX2X1 g177155(.A (n_394), .B (\cpuregs[19] [5]), .S0 (n_3216), .Y
       (n_4127));
  MX2X1 g177156(.A (n_416), .B (\cpuregs[19] [4]), .S0 (n_3216), .Y
       (n_4126));
  MX2X1 g177157(.A (n_412), .B (\cpuregs[2] [17]), .S0 (n_3218), .Y
       (n_4125));
  MX2X1 g177158(.A (n_396), .B (\cpuregs[2] [16]), .S0 (n_3218), .Y
       (n_4124));
  MX2X1 g177159(.A (n_368), .B (\cpuregs[19] [3]), .S0 (n_3216), .Y
       (n_4123));
  MX2X1 g177160(.A (n_366), .B (\cpuregs[19] [2]), .S0 (n_3216), .Y
       (n_4122));
  MX2X1 g177161(.A (n_398), .B (\cpuregs[19] [1]), .S0 (n_3216), .Y
       (n_4121));
  MX2X1 g177162(.A (n_414), .B (\cpuregs[2] [15]), .S0 (n_3218), .Y
       (n_4120));
  MX2X1 g177163(.A (n_404), .B (\cpuregs[18] [31]), .S0 (n_3217), .Y
       (n_4119));
  MX2X1 g177164(.A (n_370), .B (\cpuregs[18] [30]), .S0 (n_3217), .Y
       (n_4118));
  NAND2X1 g177165(.A (\cpuregs[2] [1]), .B (n_425), .Y (n_4117));
  AND2X1 g177166(.A (n_456), .B (\cpuregs[1] [2]), .Y (n_4116));
  AND2X1 g177167(.A (n_456), .B (\cpuregs[1] [3]), .Y (n_4115));
  NAND2X1 g177168(.A (\cpuregs[15] [7]), .B (n_462), .Y (n_4114));
  NAND2X1 g177169(.A (\cpuregs[1] [7]), .B (n_456), .Y (n_4113));
  AND2X1 g177170(.A (n_425), .B (\cpuregs[2] [14]), .Y (n_4112));
  NAND2X1 g177171(.A (\cpuregs[1] [19]), .B (n_456), .Y (n_4111));
  NAND2X1 g177172(.A (\cpuregs[1] [20]), .B (n_456), .Y (n_4110));
  NAND2X1 g177173(.A (\cpuregs[2] [22]), .B (n_425), .Y (n_4109));
  NAND2X1 g177174(.A (\cpuregs[2] [23]), .B (n_425), .Y (n_4108));
  NAND2X1 g177175(.A (\cpuregs[1] [30]), .B (n_456), .Y (n_4107));
  AND2X1 g177176(.A (n_456), .B (\cpuregs[1] [31]), .Y (n_4106));
  OR4X1 g177177(.A (\genblk2.pcpi_div_quotient_msk [26]), .B
       (\genblk2.pcpi_div_quotient_msk [24]), .C
       (\genblk2.pcpi_div_quotient_msk [23]), .D (n_3052), .Y (n_4105));
  NAND2X1 g177178(.A (n_440), .B (n_3466), .Y (n_4104));
  MX2X1 g177179(.A (n_374), .B (\cpuregs[2] [14]), .S0 (n_3218), .Y
       (n_4103));
  MX2X1 g177180(.A (n_384), .B (\cpuregs[2] [12]), .S0 (n_3218), .Y
       (n_4102));
  MX2X1 g177181(.A (n_392), .B (\cpuregs[18] [29]), .S0 (n_3217), .Y
       (n_4101));
  MX2X1 g177182(.A (n_390), .B (\cpuregs[18] [28]), .S0 (n_3217), .Y
       (n_4100));
  MX2X1 g177183(.A (n_388), .B (\cpuregs[2] [13]), .S0 (n_3218), .Y
       (n_4099));
  MX2X1 g177184(.A (n_406), .B (\cpuregs[18] [27]), .S0 (n_3217), .Y
       (n_4098));
  OAI31X1 g177185(.A0 (n_680), .A1 (n_679), .A2 (n_302), .B0 (n_3359),
       .Y (n_4097));
  OAI221X1 g177186(.A0 (n_650), .A1 (n_35), .B0 (n_683), .B1 (n_2513),
       .C0 (n_3257), .Y (n_4096));
  MX2X1 g177187(.A (n_400), .B (\cpuregs[18] [26]), .S0 (n_3217), .Y
       (n_4095));
  MX2X1 g177188(.A (n_376), .B (\cpuregs[18] [25]), .S0 (n_3217), .Y
       (n_4094));
  MX2X1 g177189(.A (n_378), .B (\cpuregs[18] [24]), .S0 (n_3217), .Y
       (n_4093));
  NOR4X1 g177190(.A (n_2593), .B (n_3129), .C (n_3128), .D (n_3127), .Y
       (n_4092));
  NOR4X1 g177191(.A (n_2594), .B (n_3126), .C (n_3106), .D (n_3125), .Y
       (n_4091));
  NOR4X1 g177192(.A (n_2587), .B (n_3120), .C (n_3165), .D (n_3118), .Y
       (n_4090));
  NOR4X1 g177193(.A (n_2591), .B (n_3108), .C (n_3107), .D (n_3105), .Y
       (n_4089));
  NOR4X1 g177194(.A (n_2592), .B (n_3094), .C (n_3093), .D (n_3092), .Y
       (n_4088));
  NOR4X1 g177195(.A (n_2590), .B (n_3088), .C (n_3087), .D (n_3086), .Y
       (n_4087));
  NOR4X1 g177196(.A (n_2588), .B (n_3083), .C (n_3082), .D (n_3081), .Y
       (n_4086));
  AOI22X1 g177197(.A0 (n_3247), .A1 (n_344), .B0 (\reg_op2[2]_9671 ),
       .B1 (n_832), .Y (n_4085));
  AOI22X1 g177198(.A0 (n_3245), .A1 (n_344), .B0 (\reg_op2[3]_9672 ),
       .B1 (n_832), .Y (n_4084));
  AOI222X1 g177199(.A0 (n_2435), .A1 (n_419), .B0 (decoded_rs2[3]), .B1
       (n_953), .C0 (n_2140), .C1 (n_3252), .Y (n_4083));
  MX2X1 g177200(.A (n_372), .B (\cpuregs[11] [9]), .S0 (n_3212), .Y
       (n_4082));
  MX2X1 g177201(.A (n_408), .B (\cpuregs[11] [10]), .S0 (n_3212), .Y
       (n_4081));
  MX2X1 g177202(.A (n_418), .B (\cpuregs[11] [8]), .S0 (n_3212), .Y
       (n_4080));
  MX2X1 g177203(.A (n_402), .B (\cpuregs[11] [11]), .S0 (n_3212), .Y
       (n_4079));
  MX2X1 g177204(.A (n_384), .B (\cpuregs[11] [12]), .S0 (n_3212), .Y
       (n_4078));
  MX2X1 g177205(.A (n_388), .B (\cpuregs[11] [13]), .S0 (n_3212), .Y
       (n_4077));
  MX2X1 g177206(.A (n_374), .B (\cpuregs[11] [14]), .S0 (n_3212), .Y
       (n_4076));
  MX2X1 g177207(.A (n_414), .B (\cpuregs[11] [15]), .S0 (n_3212), .Y
       (n_4075));
  MX2X1 g177208(.A (n_396), .B (\cpuregs[11] [16]), .S0 (n_3212), .Y
       (n_4074));
  MX2X1 g177209(.A (n_412), .B (\cpuregs[11] [17]), .S0 (n_3212), .Y
       (n_4073));
  MX2X1 g177210(.A (n_382), .B (\cpuregs[11] [18]), .S0 (n_3212), .Y
       (n_4072));
  MX2X1 g177211(.A (n_1518), .B (\cpuregs[11] [19]), .S0 (n_3212), .Y
       (n_4071));
  MX2X1 g177212(.A (n_1513), .B (\cpuregs[11] [22]), .S0 (n_3212), .Y
       (n_4070));
  MX2X1 g177213(.A (n_364), .B (\cpuregs[11] [20]), .S0 (n_3212), .Y
       (n_4069));
  MX2X1 g177214(.A (n_1515), .B (\cpuregs[11] [21]), .S0 (n_3212), .Y
       (n_4068));
  MX2X1 g177215(.A (n_380), .B (\cpuregs[11] [23]), .S0 (n_3212), .Y
       (n_4067));
  MX2X1 g177216(.A (n_378), .B (\cpuregs[11] [24]), .S0 (n_3212), .Y
       (n_4066));
  MX2X1 g177217(.A (n_376), .B (\cpuregs[11] [25]), .S0 (n_3212), .Y
       (n_4065));
  MX2X1 g177218(.A (n_400), .B (\cpuregs[11] [26]), .S0 (n_3212), .Y
       (n_4064));
  MX2X1 g177219(.A (n_406), .B (\cpuregs[11] [27]), .S0 (n_3212), .Y
       (n_4063));
  MX2X1 g177220(.A (n_390), .B (\cpuregs[11] [28]), .S0 (n_3212), .Y
       (n_4062));
  MX2X1 g177221(.A (n_392), .B (\cpuregs[11] [29]), .S0 (n_3212), .Y
       (n_4061));
  MX2X1 g177222(.A (n_370), .B (\cpuregs[11] [30]), .S0 (n_3212), .Y
       (n_4060));
  MX2X1 g177223(.A (n_398), .B (\cpuregs[13] [1]), .S0 (n_3233), .Y
       (n_4059));
  MX2X1 g177224(.A (n_366), .B (\cpuregs[13] [2]), .S0 (n_3233), .Y
       (n_4058));
  MX2X1 g177225(.A (n_368), .B (\cpuregs[13] [3]), .S0 (n_3233), .Y
       (n_4057));
  MX2X1 g177226(.A (n_416), .B (\cpuregs[13] [4]), .S0 (n_3233), .Y
       (n_4056));
  MX2X1 g177227(.A (n_394), .B (\cpuregs[13] [5]), .S0 (n_3233), .Y
       (n_4055));
  MX2X1 g177228(.A (n_362), .B (\cpuregs[13] [6]), .S0 (n_3233), .Y
       (n_4054));
  MX2X1 g177229(.A (n_386), .B (\cpuregs[13] [7]), .S0 (n_3233), .Y
       (n_4053));
  MX2X1 g177230(.A (n_418), .B (\cpuregs[13] [8]), .S0 (n_3233), .Y
       (n_4052));
  MX2X1 g177231(.A (n_372), .B (\cpuregs[13] [9]), .S0 (n_3233), .Y
       (n_4051));
  MX2X1 g177232(.A (n_408), .B (\cpuregs[13] [10]), .S0 (n_3233), .Y
       (n_4050));
  MX2X1 g177233(.A (n_402), .B (\cpuregs[13] [11]), .S0 (n_3233), .Y
       (n_4049));
  MX2X1 g177234(.A (n_384), .B (\cpuregs[13] [12]), .S0 (n_3233), .Y
       (n_4048));
  MX2X1 g177235(.A (n_388), .B (\cpuregs[13] [13]), .S0 (n_3233), .Y
       (n_4047));
  MX2X1 g177236(.A (n_414), .B (\cpuregs[13] [15]), .S0 (n_3233), .Y
       (n_4046));
  MX2X1 g177237(.A (n_374), .B (\cpuregs[13] [14]), .S0 (n_3233), .Y
       (n_4045));
  MX2X1 g177238(.A (n_396), .B (\cpuregs[13] [16]), .S0 (n_3233), .Y
       (n_4044));
  MX2X1 g177239(.A (n_412), .B (\cpuregs[13] [17]), .S0 (n_3233), .Y
       (n_4043));
  MX2X1 g177240(.A (n_382), .B (\cpuregs[13] [18]), .S0 (n_3233), .Y
       (n_4042));
  MX2X1 g177241(.A (n_1518), .B (\cpuregs[13] [19]), .S0 (n_3233), .Y
       (n_4041));
  MX2X1 g177242(.A (n_364), .B (\cpuregs[13] [20]), .S0 (n_3233), .Y
       (n_4040));
  MX2X1 g177243(.A (n_1515), .B (\cpuregs[13] [21]), .S0 (n_3233), .Y
       (n_4039));
  MX2X1 g177244(.A (n_1513), .B (\cpuregs[13] [22]), .S0 (n_3233), .Y
       (n_4038));
  MX2X1 g177245(.A (n_380), .B (\cpuregs[13] [23]), .S0 (n_3233), .Y
       (n_4037));
  MX2X1 g177246(.A (n_378), .B (\cpuregs[13] [24]), .S0 (n_3233), .Y
       (n_4036));
  MX2X1 g177248(.A (n_400), .B (\cpuregs[13] [26]), .S0 (n_3233), .Y
       (n_4035));
  MX2X1 g177249(.A (n_406), .B (\cpuregs[13] [27]), .S0 (n_3233), .Y
       (n_4034));
  MX2X1 g177250(.A (n_390), .B (\cpuregs[13] [28]), .S0 (n_3233), .Y
       (n_4033));
  MX2X1 g177251(.A (n_392), .B (\cpuregs[13] [29]), .S0 (n_3233), .Y
       (n_4032));
  MX2X1 g177252(.A (n_370), .B (\cpuregs[13] [30]), .S0 (n_3233), .Y
       (n_4031));
  MX2X1 g177253(.A (n_404), .B (\cpuregs[13] [31]), .S0 (n_3233), .Y
       (n_4030));
  MX2X1 g177254(.A (n_398), .B (\cpuregs[14] [1]), .S0 (n_3225), .Y
       (n_4029));
  MX2X1 g177255(.A (n_366), .B (\cpuregs[14] [2]), .S0 (n_3225), .Y
       (n_4028));
  MX2X1 g177256(.A (n_368), .B (\cpuregs[14] [3]), .S0 (n_3225), .Y
       (n_4027));
  MX2X1 g177257(.A (n_416), .B (\cpuregs[14] [4]), .S0 (n_3225), .Y
       (n_4026));
  MX2X1 g177258(.A (n_394), .B (\cpuregs[14] [5]), .S0 (n_3225), .Y
       (n_4025));
  MX2X1 g177259(.A (n_362), .B (\cpuregs[14] [6]), .S0 (n_3225), .Y
       (n_4024));
  MX2X1 g177260(.A (n_386), .B (\cpuregs[14] [7]), .S0 (n_3225), .Y
       (n_4023));
  MX2X1 g177261(.A (n_418), .B (\cpuregs[14] [8]), .S0 (n_3225), .Y
       (n_4022));
  MX2X1 g177262(.A (n_372), .B (\cpuregs[14] [9]), .S0 (n_3225), .Y
       (n_4021));
  MX2X1 g177263(.A (n_408), .B (\cpuregs[14] [10]), .S0 (n_3225), .Y
       (n_4020));
  MX2X1 g177264(.A (n_402), .B (\cpuregs[14] [11]), .S0 (n_3225), .Y
       (n_4019));
  MX2X1 g177265(.A (n_384), .B (\cpuregs[14] [12]), .S0 (n_3225), .Y
       (n_4018));
  MX2X1 g177266(.A (n_388), .B (\cpuregs[14] [13]), .S0 (n_3225), .Y
       (n_4017));
  MX2X1 g177267(.A (n_374), .B (\cpuregs[14] [14]), .S0 (n_3225), .Y
       (n_4016));
  MX2X1 g177268(.A (n_414), .B (\cpuregs[14] [15]), .S0 (n_3225), .Y
       (n_4015));
  MX2X1 g177269(.A (n_396), .B (\cpuregs[14] [16]), .S0 (n_3225), .Y
       (n_4014));
  MX2X1 g177270(.A (n_412), .B (\cpuregs[14] [17]), .S0 (n_3225), .Y
       (n_4013));
  MX2X1 g177271(.A (n_382), .B (\cpuregs[14] [18]), .S0 (n_3225), .Y
       (n_4012));
  MX2X1 g177272(.A (n_1518), .B (\cpuregs[14] [19]), .S0 (n_3225), .Y
       (n_4011));
  MX2X1 g177273(.A (n_364), .B (\cpuregs[14] [20]), .S0 (n_3225), .Y
       (n_4010));
  MX2X1 g177274(.A (n_1515), .B (\cpuregs[14] [21]), .S0 (n_3225), .Y
       (n_4009));
  MX2X1 g177275(.A (n_1513), .B (\cpuregs[14] [22]), .S0 (n_3225), .Y
       (n_4008));
  MX2X1 g177276(.A (n_380), .B (\cpuregs[14] [23]), .S0 (n_3225), .Y
       (n_4007));
  MX2X1 g177277(.A (n_378), .B (\cpuregs[14] [24]), .S0 (n_3225), .Y
       (n_4006));
  MX2X1 g177278(.A (n_376), .B (\cpuregs[14] [25]), .S0 (n_3225), .Y
       (n_4005));
  MX2X1 g177279(.A (n_406), .B (\cpuregs[14] [27]), .S0 (n_3225), .Y
       (n_4004));
  MX2X1 g177280(.A (n_390), .B (\cpuregs[14] [28]), .S0 (n_3225), .Y
       (n_4003));
  MX2X1 g177281(.A (n_400), .B (\cpuregs[14] [26]), .S0 (n_3225), .Y
       (n_4002));
  MX2X1 g177282(.A (n_392), .B (\cpuregs[14] [29]), .S0 (n_3225), .Y
       (n_4001));
  MX2X1 g177283(.A (n_370), .B (\cpuregs[14] [30]), .S0 (n_3225), .Y
       (n_4000));
  MX2X1 g177284(.A (n_404), .B (\cpuregs[14] [31]), .S0 (n_3225), .Y
       (n_3999));
  MX2X1 g177285(.A (n_400), .B (\cpuregs[6] [26]), .S0 (n_3215), .Y
       (n_3998));
  MX2X1 g177286(.A (n_404), .B (\cpuregs[11] [31]), .S0 (n_3212), .Y
       (n_3997));
  MX2X1 g177287(.A (n_398), .B (\cpuregs[18] [1]), .S0 (n_3217), .Y
       (n_3996));
  MX2X1 g177288(.A (n_366), .B (\cpuregs[18] [2]), .S0 (n_3217), .Y
       (n_3995));
  MX2X1 g177289(.A (n_368), .B (\cpuregs[18] [3]), .S0 (n_3217), .Y
       (n_3994));
  MX2X1 g177290(.A (n_416), .B (\cpuregs[18] [4]), .S0 (n_3217), .Y
       (n_3993));
  MX2X1 g177291(.A (n_394), .B (\cpuregs[18] [5]), .S0 (n_3217), .Y
       (n_3992));
  MX2X1 g177292(.A (n_368), .B (\cpuregs[2] [3]), .S0 (n_3218), .Y
       (n_3991));
  MX2X1 g177293(.A (n_362), .B (\cpuregs[18] [6]), .S0 (n_3217), .Y
       (n_3990));
  MX2X1 g177294(.A (n_386), .B (\cpuregs[18] [7]), .S0 (n_3217), .Y
       (n_3989));
  MX2X1 g177295(.A (n_398), .B (\cpuregs[2] [1]), .S0 (n_3218), .Y
       (n_3988));
  MX2X1 g177296(.A (n_418), .B (\cpuregs[18] [8]), .S0 (n_3217), .Y
       (n_3987));
  MX2X1 g177297(.A (n_372), .B (\cpuregs[18] [9]), .S0 (n_3217), .Y
       (n_3986));
  MX2X1 g177298(.A (n_366), .B (\cpuregs[2] [2]), .S0 (n_3218), .Y
       (n_3985));
  MX2X1 g177299(.A (n_408), .B (\cpuregs[18] [10]), .S0 (n_3217), .Y
       (n_3984));
  MX2X1 g177300(.A (n_402), .B (\cpuregs[18] [11]), .S0 (n_3217), .Y
       (n_3983));
  MX2X1 g177301(.A (n_416), .B (\cpuregs[2] [4]), .S0 (n_3218), .Y
       (n_3982));
  MX2X1 g177302(.A (n_384), .B (\cpuregs[18] [12]), .S0 (n_3217), .Y
       (n_3981));
  MX2X1 g177303(.A (n_362), .B (\cpuregs[2] [6]), .S0 (n_3218), .Y
       (n_3980));
  MX2X1 g177304(.A (n_388), .B (\cpuregs[18] [13]), .S0 (n_3217), .Y
       (n_3979));
  MX2X1 g177305(.A (n_374), .B (\cpuregs[18] [14]), .S0 (n_3217), .Y
       (n_3978));
  MX2X1 g177306(.A (n_386), .B (\cpuregs[2] [7]), .S0 (n_3218), .Y
       (n_3977));
  MX2X1 g177307(.A (n_414), .B (\cpuregs[18] [15]), .S0 (n_3217), .Y
       (n_3976));
  MX2X1 g177308(.A (n_396), .B (\cpuregs[18] [16]), .S0 (n_3217), .Y
       (n_3975));
  MX2X1 g177309(.A (n_394), .B (\cpuregs[2] [5]), .S0 (n_3218), .Y
       (n_3974));
  MX2X1 g177310(.A (n_412), .B (\cpuregs[18] [17]), .S0 (n_3217), .Y
       (n_3973));
  MX2X1 g177311(.A (n_418), .B (\cpuregs[2] [8]), .S0 (n_3218), .Y
       (n_3972));
  MX2X1 g177312(.A (n_382), .B (\cpuregs[18] [18]), .S0 (n_3217), .Y
       (n_3971));
  MX2X1 g177313(.A (n_1518), .B (\cpuregs[18] [19]), .S0 (n_3217), .Y
       (n_3970));
  MX2X1 g177314(.A (n_372), .B (\cpuregs[2] [9]), .S0 (n_3218), .Y
       (n_3969));
  MX2X1 g177315(.A (n_364), .B (\cpuregs[18] [20]), .S0 (n_3217), .Y
       (n_3968));
  MX2X1 g177316(.A (n_1515), .B (\cpuregs[18] [21]), .S0 (n_3217), .Y
       (n_3967));
  MX2X1 g177317(.A (n_408), .B (\cpuregs[2] [10]), .S0 (n_3218), .Y
       (n_3966));
  MX2X1 g177318(.A (n_1513), .B (\cpuregs[18] [22]), .S0 (n_3217), .Y
       (n_3965));
  MX2X1 g177319(.A (n_380), .B (\cpuregs[18] [23]), .S0 (n_3217), .Y
       (n_3964));
  MX2X1 g177320(.A (n_402), .B (\cpuregs[2] [11]), .S0 (n_3218), .Y
       (n_3963));
  OAI2BB1X1 g177322(.A0N (n_2569), .A1N (n_35), .B0 (n_3469), .Y
       (n_4289));
  NOR2X1 g177323(.A (n_975), .B (n_3413), .Y (n_4288));
  NAND2X1 g177325(.A (cpu_state[5]), .B (n_423), .Y (n_4287));
  MX2X1 g177494(.A (\cpuregs[7] [15]), .B (n_414), .S0 (n_510), .Y
       (n_3962));
  MX2X1 g177495(.A (n_382), .B (\cpuregs[5] [18]), .S0 (n_3221), .Y
       (n_3961));
  MX2X1 g177496(.A (n_1518), .B (\cpuregs[5] [19]), .S0 (n_3221), .Y
       (n_3960));
  MX2X1 g177497(.A (n_364), .B (\cpuregs[5] [20]), .S0 (n_3221), .Y
       (n_3959));
  MX2X1 g177498(.A (n_1515), .B (\cpuregs[5] [21]), .S0 (n_3221), .Y
       (n_3958));
  MX2X1 g177499(.A (n_380), .B (\cpuregs[5] [23]), .S0 (n_3221), .Y
       (n_3957));
  MX2X1 g177500(.A (n_1513), .B (\cpuregs[5] [22]), .S0 (n_3221), .Y
       (n_3956));
  MX2X1 g177501(.A (n_412), .B (\cpuregs[27] [17]), .S0 (n_3220), .Y
       (n_3955));
  MX2X1 g177502(.A (n_378), .B (\cpuregs[5] [24]), .S0 (n_3221), .Y
       (n_3954));
  MX2X1 g177503(.A (n_376), .B (\cpuregs[5] [25]), .S0 (n_3221), .Y
       (n_3953));
  MX2X1 g177504(.A (n_400), .B (\cpuregs[5] [26]), .S0 (n_3221), .Y
       (n_3952));
  MX2X1 g177505(.A (n_406), .B (\cpuregs[5] [27]), .S0 (n_3221), .Y
       (n_3951));
  MX2X1 g177506(.A (n_390), .B (\cpuregs[5] [28]), .S0 (n_3221), .Y
       (n_3950));
  MX2X1 g177507(.A (n_392), .B (\cpuregs[5] [29]), .S0 (n_3221), .Y
       (n_3949));
  MX2X1 g177508(.A (n_370), .B (\cpuregs[5] [30]), .S0 (n_3221), .Y
       (n_3948));
  MX2X1 g177509(.A (n_398), .B (\cpuregs[26] [1]), .S0 (n_3226), .Y
       (n_3947));
  MX2X1 g177510(.A (n_404), .B (\cpuregs[5] [31]), .S0 (n_3221), .Y
       (n_3946));
  MX2X1 g177511(.A (n_366), .B (\cpuregs[26] [2]), .S0 (n_3226), .Y
       (n_3945));
  MX2X1 g177512(.A (n_368), .B (\cpuregs[26] [3]), .S0 (n_3226), .Y
       (n_3944));
  MX2X1 g177513(.A (n_416), .B (\cpuregs[26] [4]), .S0 (n_3226), .Y
       (n_3943));
  MX2X1 g177514(.A (n_394), .B (\cpuregs[26] [5]), .S0 (n_3226), .Y
       (n_3942));
  MX2X1 g177515(.A (n_362), .B (\cpuregs[26] [6]), .S0 (n_3226), .Y
       (n_3941));
  MX2X1 g177516(.A (n_386), .B (\cpuregs[26] [7]), .S0 (n_3226), .Y
       (n_3940));
  MX2X1 g177517(.A (n_418), .B (\cpuregs[26] [8]), .S0 (n_3226), .Y
       (n_3939));
  MX2X1 g177518(.A (n_372), .B (\cpuregs[26] [9]), .S0 (n_3226), .Y
       (n_3938));
  MX2X1 g177519(.A (n_408), .B (\cpuregs[26] [10]), .S0 (n_3226), .Y
       (n_3937));
  MX2X1 g177520(.A (n_368), .B (\cpuregs[6] [3]), .S0 (n_3215), .Y
       (n_3936));
  MX2X1 g177521(.A (n_402), .B (\cpuregs[26] [11]), .S0 (n_3226), .Y
       (n_3935));
  MX2X1 g177522(.A (n_384), .B (\cpuregs[26] [12]), .S0 (n_3226), .Y
       (n_3934));
  MX2X1 g177523(.A (n_388), .B (\cpuregs[26] [13]), .S0 (n_3226), .Y
       (n_3933));
  MX2X1 g177524(.A (n_374), .B (\cpuregs[26] [14]), .S0 (n_3226), .Y
       (n_3932));
  MX2X1 g177525(.A (n_416), .B (\cpuregs[6] [4]), .S0 (n_3215), .Y
       (n_3931));
  MX2X1 g177526(.A (n_394), .B (\cpuregs[6] [5]), .S0 (n_3215), .Y
       (n_3930));
  MX2X1 g177527(.A (n_414), .B (\cpuregs[26] [15]), .S0 (n_3226), .Y
       (n_3929));
  MX2X1 g177528(.A (n_396), .B (\cpuregs[26] [16]), .S0 (n_3226), .Y
       (n_3928));
  MX2X1 g177529(.A (n_412), .B (\cpuregs[26] [17]), .S0 (n_3226), .Y
       (n_3927));
  MX2X1 g177530(.A (n_362), .B (\cpuregs[6] [6]), .S0 (n_3215), .Y
       (n_3926));
  MX2X1 g177531(.A (n_382), .B (\cpuregs[26] [18]), .S0 (n_3226), .Y
       (n_3925));
  MX2X1 g177532(.A (n_386), .B (\cpuregs[6] [7]), .S0 (n_3215), .Y
       (n_3924));
  MX2X1 g177533(.A (n_1518), .B (\cpuregs[26] [19]), .S0 (n_3226), .Y
       (n_3923));
  MX2X1 g177534(.A (n_364), .B (\cpuregs[26] [20]), .S0 (n_3226), .Y
       (n_3922));
  MX2X1 g177535(.A (n_1515), .B (\cpuregs[26] [21]), .S0 (n_3226), .Y
       (n_3921));
  MX2X1 g177536(.A (n_418), .B (\cpuregs[6] [8]), .S0 (n_3215), .Y
       (n_3920));
  MX2X1 g177537(.A (n_1513), .B (\cpuregs[26] [22]), .S0 (n_3226), .Y
       (n_3919));
  MX2X1 g177538(.A (n_380), .B (\cpuregs[26] [23]), .S0 (n_3226), .Y
       (n_3918));
  MX2X1 g177539(.A (n_372), .B (\cpuregs[6] [9]), .S0 (n_3215), .Y
       (n_3917));
  MX2X1 g177540(.A (n_378), .B (\cpuregs[26] [24]), .S0 (n_3226), .Y
       (n_3916));
  MX2X1 g177541(.A (n_408), .B (\cpuregs[6] [10]), .S0 (n_3215), .Y
       (n_3915));
  MX2X1 g177542(.A (n_376), .B (\cpuregs[26] [25]), .S0 (n_3226), .Y
       (n_3914));
  MX2X1 g177543(.A (n_402), .B (\cpuregs[6] [11]), .S0 (n_3215), .Y
       (n_3913));
  MX2X1 g177544(.A (n_400), .B (\cpuregs[26] [26]), .S0 (n_3226), .Y
       (n_3912));
  MX2X1 g177545(.A (n_406), .B (\cpuregs[26] [27]), .S0 (n_3226), .Y
       (n_3911));
  MX2X1 g177546(.A (n_390), .B (\cpuregs[26] [28]), .S0 (n_3226), .Y
       (n_3910));
  MX2X1 g177547(.A (n_384), .B (\cpuregs[6] [12]), .S0 (n_3215), .Y
       (n_3909));
  MX2X1 g177548(.A (n_392), .B (\cpuregs[26] [29]), .S0 (n_3226), .Y
       (n_3908));
  MX2X1 g177549(.A (n_370), .B (\cpuregs[26] [30]), .S0 (n_3226), .Y
       (n_3907));
  MX2X1 g177550(.A (n_388), .B (\cpuregs[6] [13]), .S0 (n_3215), .Y
       (n_3906));
  MX2X1 g177551(.A (n_404), .B (\cpuregs[26] [31]), .S0 (n_3226), .Y
       (n_3905));
  MX2X1 g177552(.A (n_374), .B (\cpuregs[6] [14]), .S0 (n_3215), .Y
       (n_3904));
  MX2X1 g177553(.A (n_366), .B (\cpuregs[27] [2]), .S0 (n_3220), .Y
       (n_3903));
  MX2X1 g177554(.A (n_414), .B (\cpuregs[6] [15]), .S0 (n_3215), .Y
       (n_3902));
  MX2X1 g177555(.A (n_416), .B (\cpuregs[27] [4]), .S0 (n_3220), .Y
       (n_3901));
  MX2X1 g177556(.A (n_394), .B (\cpuregs[27] [5]), .S0 (n_3220), .Y
       (n_3900));
  MX2X1 g177557(.A (n_412), .B (\cpuregs[6] [17]), .S0 (n_3215), .Y
       (n_3899));
  MX2X1 g177558(.A (n_362), .B (\cpuregs[27] [6]), .S0 (n_3220), .Y
       (n_3898));
  MX2X1 g177559(.A (n_386), .B (\cpuregs[27] [7]), .S0 (n_3220), .Y
       (n_3897));
  MX2X1 g177560(.A (n_382), .B (\cpuregs[6] [18]), .S0 (n_3215), .Y
       (n_3896));
  MX2X1 g177561(.A (n_418), .B (\cpuregs[27] [8]), .S0 (n_3220), .Y
       (n_3895));
  MX2X1 g177562(.A (n_408), .B (\cpuregs[27] [10]), .S0 (n_3220), .Y
       (n_3894));
  MX2X1 g177563(.A (n_396), .B (\cpuregs[6] [16]), .S0 (n_3215), .Y
       (n_3893));
  MX2X1 g177564(.A (n_402), .B (\cpuregs[27] [11]), .S0 (n_3220), .Y
       (n_3892));
  MX2X1 g177565(.A (n_1518), .B (\cpuregs[6] [19]), .S0 (n_3215), .Y
       (n_3891));
  MX2X1 g177566(.A (n_384), .B (\cpuregs[27] [12]), .S0 (n_3220), .Y
       (n_3890));
  MX2X1 g177567(.A (n_388), .B (\cpuregs[27] [13]), .S0 (n_3220), .Y
       (n_3889));
  MX2X1 g177568(.A (n_374), .B (\cpuregs[27] [14]), .S0 (n_3220), .Y
       (n_3888));
  MX2X1 g177569(.A (n_364), .B (\cpuregs[6] [20]), .S0 (n_3215), .Y
       (n_3887));
  MX2X1 g177570(.A (n_1515), .B (\cpuregs[6] [21]), .S0 (n_3215), .Y
       (n_3886));
  MX2X1 g177571(.A (n_1513), .B (\cpuregs[6] [22]), .S0 (n_3215), .Y
       (n_3885));
  MX2X1 g177572(.A (n_396), .B (\cpuregs[27] [16]), .S0 (n_3220), .Y
       (n_3884));
  MX2X1 g177573(.A (n_380), .B (\cpuregs[6] [23]), .S0 (n_3215), .Y
       (n_3883));
  MX2X1 g177574(.A (n_382), .B (\cpuregs[27] [18]), .S0 (n_3220), .Y
       (n_3882));
  MX2X1 g177575(.A (n_1518), .B (\cpuregs[27] [19]), .S0 (n_3220), .Y
       (n_3881));
  MX2X1 g177576(.A (n_364), .B (\cpuregs[27] [20]), .S0 (n_3220), .Y
       (n_3880));
  MX2X1 g177577(.A (n_378), .B (\cpuregs[6] [24]), .S0 (n_3215), .Y
       (n_3879));
  MX2X1 g177578(.A (n_1515), .B (\cpuregs[27] [21]), .S0 (n_3220), .Y
       (n_3878));
  MX2X1 g177579(.A (n_1513), .B (\cpuregs[27] [22]), .S0 (n_3220), .Y
       (n_3877));
  MX2X1 g177580(.A (n_380), .B (\cpuregs[27] [23]), .S0 (n_3220), .Y
       (n_3876));
  MX2X1 g177581(.A (n_378), .B (\cpuregs[27] [24]), .S0 (n_3220), .Y
       (n_3875));
  MX2X1 g177582(.A (n_376), .B (\cpuregs[6] [25]), .S0 (n_3215), .Y
       (n_3874));
  MX2X1 g177583(.A (n_376), .B (\cpuregs[27] [25]), .S0 (n_3220), .Y
       (n_3873));
  MX2X1 g177584(.A (n_406), .B (\cpuregs[6] [27]), .S0 (n_3215), .Y
       (n_3872));
  MX2X1 g177585(.A (n_400), .B (\cpuregs[27] [26]), .S0 (n_3220), .Y
       (n_3871));
  MX2X1 g177586(.A (n_406), .B (\cpuregs[27] [27]), .S0 (n_3220), .Y
       (n_3870));
  MX2X1 g177587(.A (n_390), .B (\cpuregs[27] [28]), .S0 (n_3220), .Y
       (n_3869));
  MX2X1 g177588(.A (n_392), .B (\cpuregs[27] [29]), .S0 (n_3220), .Y
       (n_3868));
  MX2X1 g177589(.A (n_370), .B (\cpuregs[27] [30]), .S0 (n_3220), .Y
       (n_3867));
  MX2X1 g177590(.A (n_404), .B (\cpuregs[27] [31]), .S0 (n_3220), .Y
       (n_3866));
  MX2X1 g177591(.A (n_390), .B (\cpuregs[6] [28]), .S0 (n_3215), .Y
       (n_3865));
  MX2X1 g177592(.A (n_370), .B (\cpuregs[6] [30]), .S0 (n_3215), .Y
       (n_3864));
  MX2X1 g177593(.A (n_392), .B (\cpuregs[6] [29]), .S0 (n_3215), .Y
       (n_3863));
  MX2X1 g177594(.A (n_404), .B (\cpuregs[6] [31]), .S0 (n_3215), .Y
       (n_3862));
  MX2X1 g177595(.A (n_414), .B (\cpuregs[27] [15]), .S0 (n_3220), .Y
       (n_3861));
  MX2X1 g177596(.A (n_368), .B (\cpuregs[10] [3]), .S0 (n_3229), .Y
       (n_3860));
  MX2X1 g177597(.A (n_398), .B (\cpuregs[10] [1]), .S0 (n_3229), .Y
       (n_3859));
  MX2X1 g177598(.A (n_366), .B (\cpuregs[10] [2]), .S0 (n_3229), .Y
       (n_3858));
  MX2X1 g177599(.A (n_416), .B (\cpuregs[10] [4]), .S0 (n_3229), .Y
       (n_3857));
  MX2X1 g177600(.A (n_394), .B (\cpuregs[10] [5]), .S0 (n_3229), .Y
       (n_3856));
  MX2X1 g177601(.A (n_362), .B (\cpuregs[10] [6]), .S0 (n_3229), .Y
       (n_3855));
  MX2X1 g177602(.A (n_386), .B (\cpuregs[10] [7]), .S0 (n_3229), .Y
       (n_3854));
  MX2X1 g177603(.A (n_418), .B (\cpuregs[10] [8]), .S0 (n_3229), .Y
       (n_3853));
  MX2X1 g177604(.A (n_372), .B (\cpuregs[10] [9]), .S0 (n_3229), .Y
       (n_3852));
  MX2X1 g177605(.A (n_408), .B (\cpuregs[10] [10]), .S0 (n_3229), .Y
       (n_3851));
  MX2X1 g177606(.A (n_402), .B (\cpuregs[10] [11]), .S0 (n_3229), .Y
       (n_3850));
  MX2X1 g177607(.A (n_384), .B (\cpuregs[10] [12]), .S0 (n_3229), .Y
       (n_3849));
  MX2X1 g177608(.A (n_388), .B (\cpuregs[10] [13]), .S0 (n_3229), .Y
       (n_3848));
  MX2X1 g177609(.A (n_374), .B (\cpuregs[10] [14]), .S0 (n_3229), .Y
       (n_3847));
  MX2X1 g177610(.A (n_396), .B (\cpuregs[10] [16]), .S0 (n_3229), .Y
       (n_3846));
  MX2X1 g177611(.A (n_414), .B (\cpuregs[10] [15]), .S0 (n_3229), .Y
       (n_3845));
  MX2X1 g177612(.A (n_412), .B (\cpuregs[10] [17]), .S0 (n_3229), .Y
       (n_3844));
  MX2X1 g177613(.A (n_382), .B (\cpuregs[10] [18]), .S0 (n_3229), .Y
       (n_3843));
  MX2X1 g177614(.A (n_1518), .B (\cpuregs[10] [19]), .S0 (n_3229), .Y
       (n_3842));
  MX2X1 g177615(.A (n_364), .B (\cpuregs[10] [20]), .S0 (n_3229), .Y
       (n_3841));
  MX2X1 g177616(.A (n_1513), .B (\cpuregs[10] [22]), .S0 (n_3229), .Y
       (n_3840));
  MX2X1 g177617(.A (n_1515), .B (\cpuregs[10] [21]), .S0 (n_3229), .Y
       (n_3839));
  MX2X1 g177618(.A (n_380), .B (\cpuregs[10] [23]), .S0 (n_3229), .Y
       (n_3838));
  MX2X1 g177619(.A (n_378), .B (\cpuregs[10] [24]), .S0 (n_3229), .Y
       (n_3837));
  MX2X1 g177620(.A (n_376), .B (\cpuregs[10] [25]), .S0 (n_3229), .Y
       (n_3836));
  MX2X1 g177621(.A (n_400), .B (\cpuregs[10] [26]), .S0 (n_3229), .Y
       (n_3835));
  MX2X1 g177622(.A (n_390), .B (\cpuregs[10] [28]), .S0 (n_3229), .Y
       (n_3834));
  MX2X1 g177623(.A (n_406), .B (\cpuregs[10] [27]), .S0 (n_3229), .Y
       (n_3833));
  MX2X1 g177624(.A (n_392), .B (\cpuregs[10] [29]), .S0 (n_3229), .Y
       (n_3832));
  MX2X1 g177625(.A (n_370), .B (\cpuregs[10] [30]), .S0 (n_3229), .Y
       (n_3831));
  MX2X1 g177626(.A (n_404), .B (\cpuregs[10] [31]), .S0 (n_3229), .Y
       (n_3830));
  MX2X1 g177627(.A (n_398), .B (\cpuregs[11] [1]), .S0 (n_3212), .Y
       (n_3829));
  MX2X1 g177628(.A (n_366), .B (\cpuregs[11] [2]), .S0 (n_3212), .Y
       (n_3828));
  MX2X1 g177629(.A (n_368), .B (\cpuregs[11] [3]), .S0 (n_3212), .Y
       (n_3827));
  MX2X1 g177630(.A (n_416), .B (\cpuregs[11] [4]), .S0 (n_3212), .Y
       (n_3826));
  MX2X1 g177631(.A (n_394), .B (\cpuregs[11] [5]), .S0 (n_3212), .Y
       (n_3825));
  MX2X1 g177632(.A (n_362), .B (\cpuregs[11] [6]), .S0 (n_3212), .Y
       (n_3824));
  MX2X1 g177633(.A (n_386), .B (\cpuregs[11] [7]), .S0 (n_3212), .Y
       (n_3823));
  MX2X1 g177634(.A (\cpuregs[30] [1]), .B (n_398), .S0 (n_526), .Y
       (n_3822));
  MX2X1 g177635(.A (\cpuregs[30] [2]), .B (n_366), .S0 (n_526), .Y
       (n_3821));
  MX2X1 g177636(.A (\cpuregs[30] [3]), .B (n_368), .S0 (n_526), .Y
       (n_3820));
  MX2X1 g177637(.A (\cpuregs[30] [4]), .B (n_416), .S0 (n_526), .Y
       (n_3819));
  MX2X1 g177638(.A (\cpuregs[30] [5]), .B (n_394), .S0 (n_526), .Y
       (n_3818));
  MX2X1 g177639(.A (\cpuregs[30] [6]), .B (n_362), .S0 (n_526), .Y
       (n_3817));
  MX2X1 g177640(.A (\cpuregs[30] [7]), .B (n_386), .S0 (n_526), .Y
       (n_3816));
  MX2X1 g177641(.A (\cpuregs[30] [8]), .B (n_418), .S0 (n_526), .Y
       (n_3815));
  MX2X1 g177642(.A (\cpuregs[30] [10]), .B (n_408), .S0 (n_526), .Y
       (n_3814));
  MX2X1 g177643(.A (\cpuregs[30] [11]), .B (n_402), .S0 (n_526), .Y
       (n_3813));
  MX2X1 g177644(.A (\cpuregs[30] [12]), .B (n_384), .S0 (n_526), .Y
       (n_3812));
  MX2X1 g177645(.A (\cpuregs[30] [13]), .B (n_388), .S0 (n_526), .Y
       (n_3811));
  MX2X1 g177646(.A (\cpuregs[30] [14]), .B (n_374), .S0 (n_526), .Y
       (n_3810));
  MX2X1 g177647(.A (\cpuregs[30] [9]), .B (n_372), .S0 (n_526), .Y
       (n_3809));
  MX2X1 g177648(.A (\cpuregs[30] [15]), .B (n_414), .S0 (n_526), .Y
       (n_3808));
  MX2X1 g177649(.A (\cpuregs[30] [16]), .B (n_396), .S0 (n_526), .Y
       (n_3807));
  MX2X1 g177650(.A (\cpuregs[30] [17]), .B (n_412), .S0 (n_526), .Y
       (n_3806));
  MX2X1 g177651(.A (\cpuregs[30] [18]), .B (n_382), .S0 (n_526), .Y
       (n_3805));
  MX2X1 g177652(.A (\cpuregs[30] [19]), .B (n_1518), .S0 (n_526), .Y
       (n_3804));
  MX2X1 g177653(.A (\cpuregs[30] [20]), .B (n_364), .S0 (n_526), .Y
       (n_3803));
  MX2X1 g177654(.A (\cpuregs[30] [21]), .B (n_1515), .S0 (n_526), .Y
       (n_3802));
  MX2X1 g177655(.A (\cpuregs[30] [23]), .B (n_380), .S0 (n_526), .Y
       (n_3801));
  MX2X1 g177656(.A (\cpuregs[30] [24]), .B (n_378), .S0 (n_526), .Y
       (n_3800));
  MX2X1 g177657(.A (\cpuregs[30] [22]), .B (n_1513), .S0 (n_526), .Y
       (n_3799));
  MX2X1 g177658(.A (\cpuregs[30] [26]), .B (n_400), .S0 (n_526), .Y
       (n_3798));
  MX2X1 g177659(.A (\cpuregs[30] [25]), .B (n_376), .S0 (n_526), .Y
       (n_3797));
  MX2X1 g177660(.A (\cpuregs[30] [27]), .B (n_406), .S0 (n_526), .Y
       (n_3796));
  MX2X1 g177661(.A (\cpuregs[30] [28]), .B (n_390), .S0 (n_526), .Y
       (n_3795));
  MX2X1 g177662(.A (\cpuregs[30] [30]), .B (n_370), .S0 (n_526), .Y
       (n_3794));
  MX2X1 g177663(.A (\cpuregs[30] [29]), .B (n_392), .S0 (n_526), .Y
       (n_3793));
  MX2X1 g177664(.A (\cpuregs[30] [31]), .B (n_404), .S0 (n_526), .Y
       (n_3792));
  MX2X1 g177665(.A (\cpuregs[29] [1]), .B (n_398), .S0 (n_524), .Y
       (n_3791));
  MX2X1 g177666(.A (\cpuregs[29] [2]), .B (n_366), .S0 (n_524), .Y
       (n_3790));
  MX2X1 g177667(.A (\cpuregs[29] [3]), .B (n_368), .S0 (n_524), .Y
       (n_3789));
  MX2X1 g177668(.A (\cpuregs[29] [4]), .B (n_416), .S0 (n_524), .Y
       (n_3788));
  MX2X1 g177669(.A (\cpuregs[29] [5]), .B (n_394), .S0 (n_524), .Y
       (n_3787));
  MX2X1 g177670(.A (\cpuregs[29] [6]), .B (n_362), .S0 (n_524), .Y
       (n_3786));
  MX2X1 g177671(.A (\cpuregs[29] [7]), .B (n_386), .S0 (n_524), .Y
       (n_3785));
  MX2X1 g177672(.A (\cpuregs[29] [8]), .B (n_418), .S0 (n_524), .Y
       (n_3784));
  MX2X1 g177673(.A (\cpuregs[29] [9]), .B (n_372), .S0 (n_524), .Y
       (n_3783));
  MX2X1 g177674(.A (\cpuregs[29] [10]), .B (n_408), .S0 (n_524), .Y
       (n_3782));
  MX2X1 g177675(.A (\cpuregs[29] [11]), .B (n_402), .S0 (n_524), .Y
       (n_3781));
  MX2X1 g177676(.A (\cpuregs[29] [12]), .B (n_384), .S0 (n_524), .Y
       (n_3780));
  MX2X1 g177677(.A (\cpuregs[29] [13]), .B (n_388), .S0 (n_524), .Y
       (n_3779));
  MX2X1 g177678(.A (\cpuregs[29] [14]), .B (n_374), .S0 (n_524), .Y
       (n_3778));
  MX2X1 g177679(.A (\cpuregs[29] [15]), .B (n_414), .S0 (n_524), .Y
       (n_3777));
  MX2X1 g177680(.A (\cpuregs[29] [16]), .B (n_396), .S0 (n_524), .Y
       (n_3776));
  MX2X1 g177681(.A (\cpuregs[29] [17]), .B (n_412), .S0 (n_524), .Y
       (n_3775));
  MX2X1 g177682(.A (\cpuregs[29] [18]), .B (n_382), .S0 (n_524), .Y
       (n_3774));
  MX2X1 g177683(.A (\cpuregs[29] [19]), .B (n_1518), .S0 (n_524), .Y
       (n_3773));
  MX2X1 g177684(.A (\cpuregs[29] [20]), .B (n_364), .S0 (n_524), .Y
       (n_3772));
  MX2X1 g177685(.A (\cpuregs[29] [21]), .B (n_1515), .S0 (n_524), .Y
       (n_3771));
  MX2X1 g177686(.A (\cpuregs[29] [22]), .B (n_1513), .S0 (n_524), .Y
       (n_3770));
  MX2X1 g177687(.A (\cpuregs[29] [23]), .B (n_380), .S0 (n_524), .Y
       (n_3769));
  MX2X1 g177688(.A (\cpuregs[29] [24]), .B (n_378), .S0 (n_524), .Y
       (n_3768));
  MX2X1 g177689(.A (\cpuregs[29] [25]), .B (n_376), .S0 (n_524), .Y
       (n_3767));
  MX2X1 g177690(.A (\cpuregs[29] [26]), .B (n_400), .S0 (n_524), .Y
       (n_3766));
  MX2X1 g177691(.A (\cpuregs[29] [27]), .B (n_406), .S0 (n_524), .Y
       (n_3765));
  MX2X1 g177692(.A (\cpuregs[29] [28]), .B (n_390), .S0 (n_524), .Y
       (n_3764));
  MX2X1 g177693(.A (\cpuregs[29] [29]), .B (n_392), .S0 (n_524), .Y
       (n_3763));
  MX2X1 g177694(.A (\cpuregs[29] [30]), .B (n_370), .S0 (n_524), .Y
       (n_3762));
  MX2X1 g177695(.A (\cpuregs[29] [31]), .B (n_404), .S0 (n_524), .Y
       (n_3761));
  MX2X1 g177696(.A (\cpuregs[4] [1]), .B (n_398), .S0 (n_530), .Y
       (n_3760));
  MX2X1 g177697(.A (\cpuregs[4] [2]), .B (n_366), .S0 (n_530), .Y
       (n_3759));
  MX2X1 g177698(.A (\cpuregs[4] [3]), .B (n_368), .S0 (n_530), .Y
       (n_3758));
  MX2X1 g177699(.A (\cpuregs[4] [4]), .B (n_416), .S0 (n_530), .Y
       (n_3757));
  MX2X1 g177700(.A (\cpuregs[4] [6]), .B (n_362), .S0 (n_530), .Y
       (n_3756));
  MX2X1 g177701(.A (\cpuregs[4] [5]), .B (n_394), .S0 (n_530), .Y
       (n_3755));
  MX2X1 g177702(.A (\cpuregs[4] [7]), .B (n_386), .S0 (n_530), .Y
       (n_3754));
  MX2X1 g177703(.A (\cpuregs[4] [8]), .B (n_418), .S0 (n_530), .Y
       (n_3753));
  MX2X1 g177704(.A (\cpuregs[4] [9]), .B (n_372), .S0 (n_530), .Y
       (n_3752));
  MX2X1 g177705(.A (\cpuregs[4] [10]), .B (n_408), .S0 (n_530), .Y
       (n_3751));
  MX2X1 g177706(.A (\cpuregs[4] [11]), .B (n_402), .S0 (n_530), .Y
       (n_3750));
  MX2X1 g177707(.A (\cpuregs[4] [12]), .B (n_384), .S0 (n_530), .Y
       (n_3749));
  MX2X1 g177708(.A (\cpuregs[4] [13]), .B (n_388), .S0 (n_530), .Y
       (n_3748));
  MX2X1 g177709(.A (\cpuregs[4] [14]), .B (n_374), .S0 (n_530), .Y
       (n_3747));
  MX2X1 g177710(.A (\cpuregs[4] [15]), .B (n_414), .S0 (n_530), .Y
       (n_3746));
  MX2X1 g177711(.A (\cpuregs[4] [16]), .B (n_396), .S0 (n_530), .Y
       (n_3745));
  MX2X1 g177712(.A (\cpuregs[4] [18]), .B (n_382), .S0 (n_530), .Y
       (n_3744));
  MX2X1 g177713(.A (\cpuregs[4] [17]), .B (n_412), .S0 (n_530), .Y
       (n_3743));
  MX2X1 g177714(.A (\cpuregs[4] [19]), .B (n_1518), .S0 (n_530), .Y
       (n_3742));
  MX2X1 g177715(.A (\cpuregs[4] [20]), .B (n_364), .S0 (n_530), .Y
       (n_3741));
  MX2X1 g177716(.A (\cpuregs[4] [21]), .B (n_1515), .S0 (n_530), .Y
       (n_3740));
  MX2X1 g177717(.A (\cpuregs[4] [22]), .B (n_1513), .S0 (n_530), .Y
       (n_3739));
  MX2X1 g177718(.A (\cpuregs[4] [23]), .B (n_380), .S0 (n_530), .Y
       (n_3738));
  MX2X1 g177719(.A (\cpuregs[4] [24]), .B (n_378), .S0 (n_530), .Y
       (n_3737));
  MX2X1 g177720(.A (\cpuregs[4] [25]), .B (n_376), .S0 (n_530), .Y
       (n_3736));
  MX2X1 g177721(.A (\cpuregs[4] [26]), .B (n_400), .S0 (n_530), .Y
       (n_3735));
  MX2X1 g177722(.A (\cpuregs[4] [27]), .B (n_406), .S0 (n_530), .Y
       (n_3734));
  MX2X1 g177723(.A (\cpuregs[4] [28]), .B (n_390), .S0 (n_530), .Y
       (n_3733));
  MX2X1 g177724(.A (\cpuregs[4] [29]), .B (n_392), .S0 (n_530), .Y
       (n_3732));
  MX2X1 g177725(.A (\cpuregs[4] [30]), .B (n_370), .S0 (n_530), .Y
       (n_3731));
  MX2X1 g177726(.A (\cpuregs[4] [31]), .B (n_404), .S0 (n_530), .Y
       (n_3730));
  MX2X1 g177727(.A (\cpuregs[7] [1]), .B (n_398), .S0 (n_510), .Y
       (n_3729));
  MX2X1 g177728(.A (\cpuregs[7] [3]), .B (n_368), .S0 (n_510), .Y
       (n_3728));
  MX2X1 g177729(.A (\cpuregs[7] [4]), .B (n_416), .S0 (n_510), .Y
       (n_3727));
  MX2X1 g177730(.A (\cpuregs[7] [2]), .B (n_366), .S0 (n_510), .Y
       (n_3726));
  MX2X1 g177731(.A (\cpuregs[7] [5]), .B (n_394), .S0 (n_510), .Y
       (n_3725));
  MX2X1 g177732(.A (\cpuregs[7] [6]), .B (n_362), .S0 (n_510), .Y
       (n_3724));
  MX2X1 g177733(.A (\cpuregs[7] [7]), .B (n_386), .S0 (n_510), .Y
       (n_3723));
  MX2X1 g177734(.A (\cpuregs[7] [8]), .B (n_418), .S0 (n_510), .Y
       (n_3722));
  MX2X1 g177735(.A (\cpuregs[7] [9]), .B (n_372), .S0 (n_510), .Y
       (n_3721));
  MX2X1 g177736(.A (\cpuregs[7] [10]), .B (n_408), .S0 (n_510), .Y
       (n_3720));
  MX2X1 g177737(.A (\cpuregs[7] [11]), .B (n_402), .S0 (n_510), .Y
       (n_3719));
  MX2X1 g177738(.A (\cpuregs[7] [12]), .B (n_384), .S0 (n_510), .Y
       (n_3718));
  MX2X1 g177739(.A (\cpuregs[7] [13]), .B (n_388), .S0 (n_510), .Y
       (n_3717));
  MX2X1 g177740(.A (\cpuregs[7] [14]), .B (n_374), .S0 (n_510), .Y
       (n_3716));
  MX2X1 g177741(.A (n_412), .B (\cpuregs[5] [17]), .S0 (n_3221), .Y
       (n_3715));
  MX2X1 g177742(.A (\cpuregs[7] [16]), .B (n_396), .S0 (n_510), .Y
       (n_3714));
  MX2X1 g177743(.A (\cpuregs[7] [17]), .B (n_412), .S0 (n_510), .Y
       (n_3713));
  MX2X1 g177744(.A (\cpuregs[7] [18]), .B (n_382), .S0 (n_510), .Y
       (n_3712));
  MX2X1 g177745(.A (\cpuregs[7] [19]), .B (n_1518), .S0 (n_510), .Y
       (n_3711));
  MX2X1 g177746(.A (\cpuregs[7] [20]), .B (n_364), .S0 (n_510), .Y
       (n_3710));
  MX2X1 g177747(.A (\cpuregs[7] [21]), .B (n_1515), .S0 (n_510), .Y
       (n_3709));
  MX2X1 g177748(.A (\cpuregs[7] [22]), .B (n_1513), .S0 (n_510), .Y
       (n_3708));
  MX2X1 g177749(.A (\cpuregs[7] [23]), .B (n_380), .S0 (n_510), .Y
       (n_3707));
  MX2X1 g177750(.A (\cpuregs[7] [24]), .B (n_378), .S0 (n_510), .Y
       (n_3706));
  MX2X1 g177751(.A (\cpuregs[7] [25]), .B (n_376), .S0 (n_510), .Y
       (n_3705));
  MX2X1 g177752(.A (\cpuregs[7] [26]), .B (n_400), .S0 (n_510), .Y
       (n_3704));
  MX2X1 g177753(.A (\cpuregs[7] [27]), .B (n_406), .S0 (n_510), .Y
       (n_3703));
  MX2X1 g177754(.A (\cpuregs[7] [28]), .B (n_390), .S0 (n_510), .Y
       (n_3702));
  MX2X1 g177755(.A (\cpuregs[7] [29]), .B (n_392), .S0 (n_510), .Y
       (n_3701));
  MX2X1 g177756(.A (\cpuregs[7] [30]), .B (n_370), .S0 (n_510), .Y
       (n_3700));
  MX2X1 g177757(.A (\cpuregs[7] [31]), .B (n_404), .S0 (n_510), .Y
       (n_3699));
  MX2X1 g177758(.A (\cpuregs[12] [1]), .B (n_398), .S0 (n_536), .Y
       (n_3698));
  MX2X1 g177759(.A (\cpuregs[12] [2]), .B (n_366), .S0 (n_536), .Y
       (n_3697));
  MX2X1 g177760(.A (\cpuregs[12] [3]), .B (n_368), .S0 (n_536), .Y
       (n_3696));
  MX2X1 g177761(.A (\cpuregs[12] [4]), .B (n_416), .S0 (n_536), .Y
       (n_3695));
  MX2X1 g177762(.A (\cpuregs[12] [5]), .B (n_394), .S0 (n_536), .Y
       (n_3694));
  MX2X1 g177763(.A (\cpuregs[12] [6]), .B (n_362), .S0 (n_536), .Y
       (n_3693));
  MX2X1 g177764(.A (\cpuregs[12] [8]), .B (n_418), .S0 (n_536), .Y
       (n_3692));
  MX2X1 g177765(.A (\cpuregs[12] [9]), .B (n_372), .S0 (n_536), .Y
       (n_3691));
  MX2X1 g177766(.A (\cpuregs[12] [7]), .B (n_386), .S0 (n_536), .Y
       (n_3690));
  MX2X1 g177767(.A (\cpuregs[12] [10]), .B (n_408), .S0 (n_536), .Y
       (n_3689));
  MX2X1 g177768(.A (\cpuregs[12] [11]), .B (n_402), .S0 (n_536), .Y
       (n_3688));
  MX2X1 g177769(.A (\cpuregs[12] [12]), .B (n_384), .S0 (n_536), .Y
       (n_3687));
  MX2X1 g177770(.A (\cpuregs[12] [13]), .B (n_388), .S0 (n_536), .Y
       (n_3686));
  MX2X1 g177771(.A (\cpuregs[12] [14]), .B (n_374), .S0 (n_536), .Y
       (n_3685));
  MX2X1 g177772(.A (\cpuregs[12] [15]), .B (n_414), .S0 (n_536), .Y
       (n_3684));
  MX2X1 g177773(.A (\cpuregs[12] [16]), .B (n_396), .S0 (n_536), .Y
       (n_3683));
  MX2X1 g177774(.A (\cpuregs[12] [17]), .B (n_412), .S0 (n_536), .Y
       (n_3682));
  MX2X1 g177775(.A (\cpuregs[12] [18]), .B (n_382), .S0 (n_536), .Y
       (n_3681));
  MX2X1 g177776(.A (\cpuregs[12] [19]), .B (n_1518), .S0 (n_536), .Y
       (n_3680));
  MX2X1 g177777(.A (\cpuregs[12] [20]), .B (n_364), .S0 (n_536), .Y
       (n_3679));
  MX2X1 g177778(.A (\cpuregs[12] [21]), .B (n_1515), .S0 (n_536), .Y
       (n_3678));
  MX2X1 g177779(.A (\cpuregs[12] [22]), .B (n_1513), .S0 (n_536), .Y
       (n_3677));
  MX2X1 g177780(.A (\cpuregs[12] [23]), .B (n_380), .S0 (n_536), .Y
       (n_3676));
  MX2X1 g177781(.A (\cpuregs[12] [24]), .B (n_378), .S0 (n_536), .Y
       (n_3675));
  MX2X1 g177782(.A (\cpuregs[12] [25]), .B (n_376), .S0 (n_536), .Y
       (n_3674));
  MX2X1 g177783(.A (\cpuregs[12] [26]), .B (n_400), .S0 (n_536), .Y
       (n_3673));
  MX2X1 g177784(.A (\cpuregs[12] [27]), .B (n_406), .S0 (n_536), .Y
       (n_3672));
  MX2X1 g177785(.A (\cpuregs[12] [28]), .B (n_390), .S0 (n_536), .Y
       (n_3671));
  MX2X1 g177786(.A (\cpuregs[12] [29]), .B (n_392), .S0 (n_536), .Y
       (n_3670));
  MX2X1 g177787(.A (\cpuregs[12] [30]), .B (n_370), .S0 (n_536), .Y
       (n_3669));
  MX2X1 g177788(.A (\cpuregs[12] [31]), .B (n_404), .S0 (n_536), .Y
       (n_3668));
  MX2X1 g177789(.A (\cpuregs[15] [2]), .B (n_366), .S0 (n_512), .Y
       (n_3667));
  MX2X1 g177790(.A (\cpuregs[15] [1]), .B (n_398), .S0 (n_512), .Y
       (n_3666));
  MX2X1 g177791(.A (\cpuregs[15] [3]), .B (n_368), .S0 (n_512), .Y
       (n_3665));
  MX2X1 g177792(.A (\cpuregs[15] [4]), .B (n_416), .S0 (n_512), .Y
       (n_3664));
  MX2X1 g177793(.A (\cpuregs[15] [5]), .B (n_394), .S0 (n_512), .Y
       (n_3663));
  MX2X1 g177794(.A (\cpuregs[15] [6]), .B (n_362), .S0 (n_512), .Y
       (n_3662));
  MX2X1 g177795(.A (\cpuregs[15] [7]), .B (n_386), .S0 (n_512), .Y
       (n_3661));
  MX2X1 g177796(.A (\cpuregs[15] [8]), .B (n_418), .S0 (n_512), .Y
       (n_3660));
  MX2X1 g177797(.A (\cpuregs[15] [9]), .B (n_372), .S0 (n_512), .Y
       (n_3659));
  MX2X1 g177798(.A (\cpuregs[15] [10]), .B (n_408), .S0 (n_512), .Y
       (n_3658));
  MX2X1 g177799(.A (\cpuregs[15] [11]), .B (n_402), .S0 (n_512), .Y
       (n_3657));
  MX2X1 g177800(.A (\cpuregs[15] [12]), .B (n_384), .S0 (n_512), .Y
       (n_3656));
  MX2X1 g177801(.A (\cpuregs[15] [13]), .B (n_388), .S0 (n_512), .Y
       (n_3655));
  MX2X1 g177802(.A (\cpuregs[15] [14]), .B (n_374), .S0 (n_512), .Y
       (n_3654));
  MX2X1 g177803(.A (\cpuregs[15] [15]), .B (n_414), .S0 (n_512), .Y
       (n_3653));
  MX2X1 g177804(.A (\cpuregs[15] [16]), .B (n_396), .S0 (n_512), .Y
       (n_3652));
  MX2X1 g177805(.A (\cpuregs[15] [17]), .B (n_412), .S0 (n_512), .Y
       (n_3651));
  MX2X1 g177806(.A (\cpuregs[15] [18]), .B (n_382), .S0 (n_512), .Y
       (n_3650));
  MX2X1 g177807(.A (\cpuregs[15] [19]), .B (n_1518), .S0 (n_512), .Y
       (n_3649));
  MX2X1 g177808(.A (\cpuregs[15] [20]), .B (n_364), .S0 (n_512), .Y
       (n_3648));
  MX2X1 g177809(.A (\cpuregs[15] [21]), .B (n_1515), .S0 (n_512), .Y
       (n_3647));
  MX2X1 g177810(.A (\cpuregs[15] [22]), .B (n_1513), .S0 (n_512), .Y
       (n_3646));
  MX2X1 g177811(.A (\cpuregs[15] [23]), .B (n_380), .S0 (n_512), .Y
       (n_3645));
  MX2X1 g177812(.A (\cpuregs[15] [24]), .B (n_378), .S0 (n_512), .Y
       (n_3644));
  MX2X1 g177813(.A (\cpuregs[15] [25]), .B (n_376), .S0 (n_512), .Y
       (n_3643));
  MX2X1 g177814(.A (\cpuregs[15] [26]), .B (n_400), .S0 (n_512), .Y
       (n_3642));
  MX2X1 g177815(.A (\cpuregs[15] [27]), .B (n_406), .S0 (n_512), .Y
       (n_3641));
  MX2X1 g177816(.A (\cpuregs[15] [28]), .B (n_390), .S0 (n_512), .Y
       (n_3640));
  MX2X1 g177817(.A (\cpuregs[15] [29]), .B (n_392), .S0 (n_512), .Y
       (n_3639));
  MX2X1 g177818(.A (\cpuregs[15] [30]), .B (n_370), .S0 (n_512), .Y
       (n_3638));
  MX2X1 g177819(.A (\cpuregs[15] [31]), .B (n_404), .S0 (n_512), .Y
       (n_3637));
  MX2X1 g177820(.A (\cpuregs[20] [1]), .B (n_398), .S0 (n_532), .Y
       (n_3636));
  MX2X1 g177821(.A (\cpuregs[20] [2]), .B (n_366), .S0 (n_532), .Y
       (n_3635));
  MX2X1 g177822(.A (\cpuregs[20] [3]), .B (n_368), .S0 (n_532), .Y
       (n_3634));
  MX2X1 g177823(.A (\cpuregs[20] [4]), .B (n_416), .S0 (n_532), .Y
       (n_3633));
  MX2X1 g177824(.A (\cpuregs[20] [5]), .B (n_394), .S0 (n_532), .Y
       (n_3632));
  MX2X1 g177825(.A (\cpuregs[20] [6]), .B (n_362), .S0 (n_532), .Y
       (n_3631));
  MX2X1 g177826(.A (\cpuregs[20] [7]), .B (n_386), .S0 (n_532), .Y
       (n_3630));
  MX2X1 g177827(.A (\cpuregs[20] [8]), .B (n_418), .S0 (n_532), .Y
       (n_3629));
  MX2X1 g177828(.A (\cpuregs[20] [9]), .B (n_372), .S0 (n_532), .Y
       (n_3628));
  MX2X1 g177829(.A (\cpuregs[20] [10]), .B (n_408), .S0 (n_532), .Y
       (n_3627));
  MX2X1 g177830(.A (\cpuregs[20] [11]), .B (n_402), .S0 (n_532), .Y
       (n_3626));
  MX2X1 g177831(.A (\cpuregs[20] [12]), .B (n_384), .S0 (n_532), .Y
       (n_3625));
  MX2X1 g177832(.A (\cpuregs[20] [13]), .B (n_388), .S0 (n_532), .Y
       (n_3624));
  MX2X1 g177833(.A (\cpuregs[20] [14]), .B (n_374), .S0 (n_532), .Y
       (n_3623));
  MX2X1 g177834(.A (\cpuregs[20] [15]), .B (n_414), .S0 (n_532), .Y
       (n_3622));
  MX2X1 g177835(.A (\cpuregs[20] [16]), .B (n_396), .S0 (n_532), .Y
       (n_3621));
  MX2X1 g177836(.A (\cpuregs[20] [17]), .B (n_412), .S0 (n_532), .Y
       (n_3620));
  MX2X1 g177837(.A (\cpuregs[20] [18]), .B (n_382), .S0 (n_532), .Y
       (n_3619));
  MX2X1 g177838(.A (\cpuregs[20] [19]), .B (n_1518), .S0 (n_532), .Y
       (n_3618));
  MX2X1 g177839(.A (\cpuregs[20] [20]), .B (n_364), .S0 (n_532), .Y
       (n_3617));
  MX2X1 g177840(.A (\cpuregs[20] [21]), .B (n_1515), .S0 (n_532), .Y
       (n_3616));
  MX2X1 g177841(.A (\cpuregs[20] [22]), .B (n_1513), .S0 (n_532), .Y
       (n_3615));
  MX2X1 g177842(.A (\cpuregs[20] [23]), .B (n_380), .S0 (n_532), .Y
       (n_3614));
  MX2X1 g177843(.A (\cpuregs[20] [24]), .B (n_378), .S0 (n_532), .Y
       (n_3613));
  MX2X1 g177844(.A (\cpuregs[20] [25]), .B (n_376), .S0 (n_532), .Y
       (n_3612));
  MX2X1 g177845(.A (\cpuregs[20] [26]), .B (n_400), .S0 (n_532), .Y
       (n_3611));
  MX2X1 g177846(.A (\cpuregs[20] [27]), .B (n_406), .S0 (n_532), .Y
       (n_3610));
  MX2X1 g177847(.A (\cpuregs[20] [28]), .B (n_390), .S0 (n_532), .Y
       (n_3609));
  MX2X1 g177848(.A (\cpuregs[20] [29]), .B (n_392), .S0 (n_532), .Y
       (n_3608));
  MX2X1 g177849(.A (\cpuregs[20] [30]), .B (n_370), .S0 (n_532), .Y
       (n_3607));
  MX2X1 g177850(.A (\cpuregs[20] [31]), .B (n_404), .S0 (n_532), .Y
       (n_3606));
  MX2X1 g177851(.A (\cpuregs[23] [1]), .B (n_398), .S0 (n_518), .Y
       (n_3605));
  MX2X1 g177852(.A (\cpuregs[23] [2]), .B (n_366), .S0 (n_518), .Y
       (n_3604));
  MX2X1 g177853(.A (\cpuregs[23] [3]), .B (n_368), .S0 (n_518), .Y
       (n_3603));
  MX2X1 g177854(.A (\cpuregs[23] [4]), .B (n_416), .S0 (n_518), .Y
       (n_3602));
  MX2X1 g177855(.A (\cpuregs[23] [5]), .B (n_394), .S0 (n_518), .Y
       (n_3601));
  MX2X1 g177856(.A (\cpuregs[23] [6]), .B (n_362), .S0 (n_518), .Y
       (n_3600));
  MX2X1 g177857(.A (\cpuregs[23] [7]), .B (n_386), .S0 (n_518), .Y
       (n_3599));
  MX2X1 g177858(.A (\cpuregs[23] [8]), .B (n_418), .S0 (n_518), .Y
       (n_3598));
  MX2X1 g177859(.A (\cpuregs[23] [9]), .B (n_372), .S0 (n_518), .Y
       (n_3597));
  MX2X1 g177860(.A (\cpuregs[23] [10]), .B (n_408), .S0 (n_518), .Y
       (n_3596));
  MX2X1 g177861(.A (\cpuregs[23] [11]), .B (n_402), .S0 (n_518), .Y
       (n_3595));
  MX2X1 g177862(.A (\cpuregs[23] [12]), .B (n_384), .S0 (n_518), .Y
       (n_3594));
  MX2X1 g177863(.A (\cpuregs[23] [13]), .B (n_388), .S0 (n_518), .Y
       (n_3593));
  MX2X1 g177864(.A (\cpuregs[23] [14]), .B (n_374), .S0 (n_518), .Y
       (n_3592));
  MX2X1 g177865(.A (\cpuregs[23] [15]), .B (n_414), .S0 (n_518), .Y
       (n_3591));
  MX2X1 g177866(.A (\cpuregs[23] [16]), .B (n_396), .S0 (n_518), .Y
       (n_3590));
  MX2X1 g177867(.A (\cpuregs[23] [17]), .B (n_412), .S0 (n_518), .Y
       (n_3589));
  MX2X1 g177868(.A (\cpuregs[23] [18]), .B (n_382), .S0 (n_518), .Y
       (n_3588));
  MX2X1 g177869(.A (\cpuregs[23] [19]), .B (n_1518), .S0 (n_518), .Y
       (n_3587));
  MX2X1 g177870(.A (\cpuregs[23] [20]), .B (n_364), .S0 (n_518), .Y
       (n_3586));
  MX2X1 g177871(.A (\cpuregs[23] [21]), .B (n_1515), .S0 (n_518), .Y
       (n_3585));
  MX2X1 g177872(.A (\cpuregs[23] [22]), .B (n_1513), .S0 (n_518), .Y
       (n_3584));
  MX2X1 g177873(.A (\cpuregs[23] [23]), .B (n_380), .S0 (n_518), .Y
       (n_3583));
  MX2X1 g177874(.A (\cpuregs[23] [24]), .B (n_378), .S0 (n_518), .Y
       (n_3582));
  MX2X1 g177875(.A (\cpuregs[23] [25]), .B (n_376), .S0 (n_518), .Y
       (n_3581));
  MX2X1 g177876(.A (\cpuregs[23] [26]), .B (n_400), .S0 (n_518), .Y
       (n_3580));
  MX2X1 g177877(.A (\cpuregs[23] [27]), .B (n_406), .S0 (n_518), .Y
       (n_3579));
  MX2X1 g177878(.A (\cpuregs[23] [28]), .B (n_390), .S0 (n_518), .Y
       (n_3578));
  MX2X1 g177879(.A (\cpuregs[23] [29]), .B (n_392), .S0 (n_518), .Y
       (n_3577));
  MX2X1 g177880(.A (\cpuregs[23] [30]), .B (n_370), .S0 (n_518), .Y
       (n_3576));
  MX2X1 g177881(.A (\cpuregs[23] [31]), .B (n_404), .S0 (n_518), .Y
       (n_3575));
  MX2X1 g177882(.A (n_358), .B (\cpuregs[13] [0]), .S0 (n_3233), .Y
       (n_3574));
  MX2X1 g177883(.A (n_358), .B (\cpuregs[14] [0]), .S0 (n_3225), .Y
       (n_3573));
  MX2X1 g177884(.A (n_358), .B (\cpuregs[18] [0]), .S0 (n_3217), .Y
       (n_3572));
  MX2X1 g177885(.A (n_358), .B (\cpuregs[2] [0]), .S0 (n_3218), .Y
       (n_3571));
  MX2X1 g177886(.A (n_358), .B (\cpuregs[19] [0]), .S0 (n_3216), .Y
       (n_3570));
  MX2X1 g177887(.A (\cpuregs[3] [0]), .B (n_358), .S0 (n_697), .Y
       (n_3569));
  MX2X1 g177888(.A (n_358), .B (\cpuregs[21] [0]), .S0 (n_3214), .Y
       (n_3568));
  MX2X1 g177889(.A (n_358), .B (\cpuregs[22] [0]), .S0 (n_3213), .Y
       (n_3567));
  MX2X1 g177890(.A (n_358), .B (\cpuregs[5] [0]), .S0 (n_3221), .Y
       (n_3566));
  MX2X1 g177891(.A (n_358), .B (\cpuregs[26] [0]), .S0 (n_3226), .Y
       (n_3565));
  MX2X1 g177892(.A (n_358), .B (\cpuregs[6] [0]), .S0 (n_3215), .Y
       (n_3564));
  MX2X1 g177893(.A (n_358), .B (\cpuregs[27] [0]), .S0 (n_3220), .Y
       (n_3563));
  MX2X1 g177894(.A (n_358), .B (\cpuregs[10] [0]), .S0 (n_3229), .Y
       (n_3562));
  MX2X1 g177895(.A (n_358), .B (\cpuregs[11] [0]), .S0 (n_3212), .Y
       (n_3561));
  MX2X1 g177896(.A (\cpuregs[28] [1]), .B (n_398), .S0 (n_534), .Y
       (n_3560));
  MX2X1 g177897(.A (\cpuregs[28] [2]), .B (n_366), .S0 (n_534), .Y
       (n_3559));
  MX2X1 g177898(.A (\cpuregs[28] [3]), .B (n_368), .S0 (n_534), .Y
       (n_3558));
  MX2X1 g177899(.A (\cpuregs[28] [4]), .B (n_416), .S0 (n_534), .Y
       (n_3557));
  MX2X1 g177900(.A (\cpuregs[28] [5]), .B (n_394), .S0 (n_534), .Y
       (n_3556));
  MX2X1 g177901(.A (\cpuregs[28] [6]), .B (n_362), .S0 (n_534), .Y
       (n_3555));
  MX2X1 g177902(.A (\cpuregs[28] [7]), .B (n_386), .S0 (n_534), .Y
       (n_3554));
  MX2X1 g177903(.A (\cpuregs[28] [8]), .B (n_418), .S0 (n_534), .Y
       (n_3553));
  MX2X1 g177904(.A (\cpuregs[28] [9]), .B (n_372), .S0 (n_534), .Y
       (n_3552));
  MX2X1 g177905(.A (\cpuregs[28] [10]), .B (n_408), .S0 (n_534), .Y
       (n_3551));
  MX2X1 g177906(.A (\cpuregs[28] [11]), .B (n_402), .S0 (n_534), .Y
       (n_3550));
  MX2X1 g177907(.A (\cpuregs[28] [12]), .B (n_384), .S0 (n_534), .Y
       (n_3549));
  MX2X1 g177908(.A (\cpuregs[28] [13]), .B (n_388), .S0 (n_534), .Y
       (n_3548));
  MX2X1 g177909(.A (\cpuregs[28] [14]), .B (n_374), .S0 (n_534), .Y
       (n_3547));
  MX2X1 g177910(.A (\cpuregs[28] [15]), .B (n_414), .S0 (n_534), .Y
       (n_3546));
  MX2X1 g177911(.A (\cpuregs[28] [16]), .B (n_396), .S0 (n_534), .Y
       (n_3545));
  MX2X1 g177912(.A (\cpuregs[28] [17]), .B (n_412), .S0 (n_534), .Y
       (n_3544));
  MX2X1 g177913(.A (\cpuregs[28] [18]), .B (n_382), .S0 (n_534), .Y
       (n_3543));
  MX2X1 g177914(.A (\cpuregs[28] [19]), .B (n_1518), .S0 (n_534), .Y
       (n_3542));
  MX2X1 g177915(.A (\cpuregs[28] [20]), .B (n_364), .S0 (n_534), .Y
       (n_3541));
  MX2X1 g177916(.A (\cpuregs[28] [21]), .B (n_1515), .S0 (n_534), .Y
       (n_3540));
  MX2X1 g177917(.A (\cpuregs[28] [22]), .B (n_1513), .S0 (n_534), .Y
       (n_3539));
  MX2X1 g177918(.A (\cpuregs[28] [23]), .B (n_380), .S0 (n_534), .Y
       (n_3538));
  MX2X1 g177919(.A (\cpuregs[28] [24]), .B (n_378), .S0 (n_534), .Y
       (n_3537));
  MX2X1 g177920(.A (\cpuregs[28] [25]), .B (n_376), .S0 (n_534), .Y
       (n_3536));
  MX2X1 g177921(.A (\cpuregs[28] [26]), .B (n_400), .S0 (n_534), .Y
       (n_3535));
  MX2X1 g177922(.A (\cpuregs[28] [27]), .B (n_406), .S0 (n_534), .Y
       (n_3534));
  MX2X1 g177923(.A (\cpuregs[28] [28]), .B (n_390), .S0 (n_534), .Y
       (n_3533));
  MX2X1 g177924(.A (\cpuregs[28] [29]), .B (n_392), .S0 (n_534), .Y
       (n_3532));
  MX2X1 g177925(.A (\cpuregs[28] [30]), .B (n_370), .S0 (n_534), .Y
       (n_3531));
  MX2X1 g177926(.A (\cpuregs[28] [31]), .B (n_404), .S0 (n_534), .Y
       (n_3530));
  MX2X1 g177927(.A (\cpuregs[31] [1]), .B (n_398), .S0 (n_528), .Y
       (n_3529));
  MX2X1 g177928(.A (\cpuregs[31] [2]), .B (n_366), .S0 (n_528), .Y
       (n_3528));
  MX2X1 g177929(.A (\cpuregs[31] [3]), .B (n_368), .S0 (n_528), .Y
       (n_3527));
  MX2X1 g177930(.A (\cpuregs[31] [4]), .B (n_416), .S0 (n_528), .Y
       (n_3526));
  MX2X1 g177931(.A (\cpuregs[31] [5]), .B (n_394), .S0 (n_528), .Y
       (n_3525));
  MX2X1 g177932(.A (\cpuregs[31] [6]), .B (n_362), .S0 (n_528), .Y
       (n_3524));
  MX2X1 g177933(.A (\cpuregs[31] [7]), .B (n_386), .S0 (n_528), .Y
       (n_3523));
  MX2X1 g177934(.A (\cpuregs[31] [8]), .B (n_418), .S0 (n_528), .Y
       (n_3522));
  MX2X1 g177935(.A (\cpuregs[31] [9]), .B (n_372), .S0 (n_528), .Y
       (n_3521));
  MX2X1 g177936(.A (\cpuregs[31] [10]), .B (n_408), .S0 (n_528), .Y
       (n_3520));
  MX2X1 g177937(.A (\cpuregs[31] [11]), .B (n_402), .S0 (n_528), .Y
       (n_3519));
  MX2X1 g177938(.A (\cpuregs[31] [12]), .B (n_384), .S0 (n_528), .Y
       (n_3518));
  MX2X1 g177939(.A (\cpuregs[31] [13]), .B (n_388), .S0 (n_528), .Y
       (n_3517));
  MX2X1 g177940(.A (\cpuregs[31] [14]), .B (n_374), .S0 (n_528), .Y
       (n_3516));
  MX2X1 g177941(.A (\cpuregs[31] [15]), .B (n_414), .S0 (n_528), .Y
       (n_3515));
  MX2X1 g177942(.A (\cpuregs[31] [16]), .B (n_396), .S0 (n_528), .Y
       (n_3514));
  MX2X1 g177943(.A (\cpuregs[31] [17]), .B (n_412), .S0 (n_528), .Y
       (n_3513));
  MX2X1 g177944(.A (\cpuregs[31] [18]), .B (n_382), .S0 (n_528), .Y
       (n_3512));
  MX2X1 g177945(.A (\cpuregs[31] [19]), .B (n_1518), .S0 (n_528), .Y
       (n_3511));
  MX2X1 g177946(.A (\cpuregs[31] [21]), .B (n_1515), .S0 (n_528), .Y
       (n_3510));
  MX2X1 g177947(.A (\cpuregs[31] [20]), .B (n_364), .S0 (n_528), .Y
       (n_3509));
  MX2X1 g177948(.A (\cpuregs[31] [22]), .B (n_1513), .S0 (n_528), .Y
       (n_3508));
  MX2X1 g177949(.A (\cpuregs[31] [23]), .B (n_380), .S0 (n_528), .Y
       (n_3507));
  MX2X1 g177950(.A (\cpuregs[31] [24]), .B (n_378), .S0 (n_528), .Y
       (n_3506));
  MX2X1 g177951(.A (\cpuregs[31] [25]), .B (n_376), .S0 (n_528), .Y
       (n_3505));
  MX2X1 g177952(.A (\cpuregs[31] [26]), .B (n_400), .S0 (n_528), .Y
       (n_3504));
  MX2X1 g177953(.A (\cpuregs[31] [27]), .B (n_406), .S0 (n_528), .Y
       (n_3503));
  MX2X1 g177954(.A (\cpuregs[31] [28]), .B (n_390), .S0 (n_528), .Y
       (n_3502));
  MX2X1 g177955(.A (\cpuregs[31] [30]), .B (n_370), .S0 (n_528), .Y
       (n_3501));
  MX2X1 g177956(.A (\cpuregs[31] [29]), .B (n_392), .S0 (n_528), .Y
       (n_3500));
  MX2X1 g177957(.A (\cpuregs[31] [31]), .B (n_404), .S0 (n_528), .Y
       (n_3499));
  MX2X1 g177958(.A (\cpuregs[30] [0]), .B (n_358), .S0 (n_526), .Y
       (n_3498));
  MX2X1 g177959(.A (\cpuregs[29] [0]), .B (n_358), .S0 (n_524), .Y
       (n_3497));
  MX2X1 g177960(.A (\cpuregs[4] [0]), .B (n_358), .S0 (n_530), .Y
       (n_3496));
  AOI211XL g177961(.A0 (is_alu_reg_imm), .A1 (n_953), .B0 (n_2612), .C0
       (n_3414), .Y (n_3495));
  MX2X1 g177962(.A (\cpuregs[7] [0]), .B (n_358), .S0 (n_510), .Y
       (n_3494));
  MX2X1 g177963(.A (\cpuregs[12] [0]), .B (n_358), .S0 (n_536), .Y
       (n_3493));
  MX2X1 g177964(.A (\cpuregs[15] [0]), .B (n_358), .S0 (n_512), .Y
       (n_3492));
  MX2X1 g177965(.A (\cpuregs[20] [0]), .B (n_358), .S0 (n_532), .Y
       (n_3491));
  MX2X1 g177966(.A (\cpuregs[23] [0]), .B (n_358), .S0 (n_518), .Y
       (n_3490));
  AOI221X1 g177967(.A0 (\cpuregs[27] [8]), .A1 (n_2525), .B0
       (\cpuregs[30] [8]), .B1 (n_2523), .C0 (n_3130), .Y (n_3489));
  AOI221X1 g177968(.A0 (\cpuregs[29] [9]), .A1 (n_2524), .B0
       (\cpuregs[28] [9]), .B1 (n_2491), .C0 (n_3121), .Y (n_3488));
  AOI221X1 g177969(.A0 (\cpuregs[26] [11]), .A1 (n_2493), .B0
       (\cpuregs[30] [11]), .B1 (n_2523), .C0 (n_3116), .Y (n_3487));
  AOI221X1 g177970(.A0 (\cpuregs[26] [12]), .A1 (n_2493), .B0
       (\cpuregs[28] [12]), .B1 (n_2491), .C0 (n_3133), .Y (n_3486));
  AOI221X1 g177971(.A0 (\cpuregs[18] [13]), .A1 (n_2519), .B0
       (\cpuregs[15] [13]), .B1 (n_2504), .C0 (n_3114), .Y (n_3485));
  AOI221X1 g177972(.A0 (\cpuregs[24] [14]), .A1 (n_2490), .B0
       (\cpuregs[28] [14]), .B1 (n_2491), .C0 (n_3112), .Y (n_3484));
  AOI221X1 g177973(.A0 (\cpuregs[29] [15]), .A1 (n_2524), .B0
       (\cpuregs[28] [15]), .B1 (n_2491), .C0 (n_3110), .Y (n_3483));
  AOI221X1 g177974(.A0 (\cpuregs[20] [16]), .A1 (n_2522), .B0
       (\cpuregs[15] [16]), .B1 (n_2504), .C0 (n_3109), .Y (n_3482));
  AOI221X1 g177975(.A0 (\cpuregs[26] [18]), .A1 (n_2493), .B0
       (\cpuregs[28] [18]), .B1 (n_2491), .C0 (n_3103), .Y (n_3481));
  AOI221X1 g177976(.A0 (\cpuregs[26] [19]), .A1 (n_2493), .B0
       (\cpuregs[30] [19]), .B1 (n_2523), .C0 (n_3101), .Y (n_3480));
  AOI221X1 g177977(.A0 (\cpuregs[22] [20]), .A1 (n_2518), .B0
       (\cpuregs[15] [20]), .B1 (n_2504), .C0 (n_3099), .Y (n_3479));
  AOI221X1 g177978(.A0 (\cpuregs[26] [21]), .A1 (n_2493), .B0
       (\cpuregs[30] [21]), .B1 (n_2523), .C0 (n_3097), .Y (n_3478));
  AOI221X1 g177979(.A0 (\cpuregs[26] [22]), .A1 (n_2493), .B0
       (\cpuregs[28] [22]), .B1 (n_2491), .C0 (n_3095), .Y (n_3477));
  AOI221X1 g177980(.A0 (\cpuregs[27] [25]), .A1 (n_2525), .B0
       (\cpuregs[30] [25]), .B1 (n_2523), .C0 (n_3089), .Y (n_3476));
  AOI221X1 g177981(.A0 (\cpuregs[27] [27]), .A1 (n_2525), .B0
       (\cpuregs[30] [27]), .B1 (n_2523), .C0 (n_3084), .Y (n_3475));
  AOI221X1 g177982(.A0 (\cpuregs[16] [30]), .A1 (n_2502), .B0
       (\cpuregs[17] [30]), .B1 (n_2527), .C0 (n_3079), .Y (n_3474));
  AOI221X1 g177983(.A0 (\cpuregs[24] [31]), .A1 (n_2490), .B0
       (\cpuregs[28] [31]), .B1 (n_2491), .C0 (n_3077), .Y (n_3473));
  MX2X1 g177984(.A (\cpuregs[28] [0]), .B (n_358), .S0 (n_534), .Y
       (n_3472));
  MX2X1 g177985(.A (\cpuregs[31] [0]), .B (n_358), .S0 (n_528), .Y
       (n_3471));
  OAI222X1 g177986(.A0 (n_611), .A1 (n_2392), .B0 (n_3246), .B1
       (n_2442), .C0 (n_646), .C1 (n_969), .Y (n_3470));
  INVX1 g177989(.A (n_3467), .Y (n_3468));
  MX2X1 g177994(.A (n_400), .B (\cpuregs[9] [26]), .S0 (n_3040), .Y
       (n_3433));
  MX2X1 g177995(.A (n_376), .B (\cpuregs[9] [25]), .S0 (n_3040), .Y
       (n_3432));
  MX2X1 g177996(.A (n_378), .B (\cpuregs[9] [24]), .S0 (n_3040), .Y
       (n_3431));
  AND2X1 g177997(.A (n_3251), .B (n_983), .Y (n_3430));
  NAND2X1 g177998(.A (n_2602), .B (n_3170), .Y (n_3429));
  MX2X1 g177999(.A (n_1515), .B (\cpuregs[9] [21]), .S0 (n_3040), .Y
       (n_3428));
  MX2X1 g178000(.A (n_380), .B (\cpuregs[9] [23]), .S0 (n_3040), .Y
       (n_3427));
  MX2X1 g178001(.A (n_1513), .B (\cpuregs[9] [22]), .S0 (n_3040), .Y
       (n_3426));
  OAI2BB1X1 g178002(.A0N (n_6534), .A1N (n_3051), .B0 (n_6541), .Y
       (n_3425));
  NAND2X1 g178003(.A (n_3044), .B (n_3075), .Y (n_3424));
  MX2X1 g178004(.A (n_412), .B (\cpuregs[9] [17]), .S0 (n_3040), .Y
       (n_3423));
  MX2X1 g178005(.A (n_364), .B (\cpuregs[9] [20]), .S0 (n_3040), .Y
       (n_3422));
  MX2X1 g178006(.A (n_1518), .B (\cpuregs[9] [19]), .S0 (n_3040), .Y
       (n_3421));
  MX2X1 g178007(.A (n_382), .B (\cpuregs[9] [18]), .S0 (n_3040), .Y
       (n_3420));
  AND2X1 g178008(.A (n_3249), .B (n_2424), .Y (n_3419));
  OAI31X1 g178009(.A0 (n_2997), .A1 (n_2610), .A2 (n_1590), .B0
       (n_2505), .Y (n_3418));
  MX2X1 g178010(.A (n_414), .B (\cpuregs[9] [15]), .S0 (n_3040), .Y
       (n_3417));
  MX2X1 g178011(.A (n_396), .B (\cpuregs[9] [16]), .S0 (n_3040), .Y
       (n_3416));
  OAI21X1 g178012(.A0 (n_14), .A1 (n_3071), .B0 (n_2140), .Y (n_3415));
  OAI2BB1X1 g178013(.A0N (n_2599), .A1N (n_1588), .B0 (n_3173), .Y
       (n_3414));
  NOR3BX1 g178014(.AN (n_1351), .B (n_849), .C (n_303), .Y (n_3413));
  OAI211X1 g178015(.A0 (n_2423), .A1 (n_2996), .B0 (n_2322), .C0
       (n_1588), .Y (n_3412));
  OAI2BB1X1 g178016(.A0N (cpu_state[3]), .A1N (n_115), .B0 (n_3168), .Y
       (n_3411));
  MX2X1 g178017(.A (n_374), .B (\cpuregs[9] [14]), .S0 (n_3040), .Y
       (n_3410));
  MX2X1 g178018(.A (n_398), .B (\cpuregs[9] [1]), .S0 (n_3040), .Y
       (n_3409));
  MX2X1 g178019(.A (n_366), .B (\cpuregs[9] [2]), .S0 (n_3040), .Y
       (n_3408));
  MX2X1 g178020(.A (n_416), .B (\cpuregs[9] [4]), .S0 (n_3040), .Y
       (n_3407));
  MX2X1 g178021(.A (n_368), .B (\cpuregs[9] [3]), .S0 (n_3040), .Y
       (n_3406));
  MX2X1 g178022(.A (n_394), .B (\cpuregs[9] [5]), .S0 (n_3040), .Y
       (n_3405));
  MX2X1 g178023(.A (n_362), .B (\cpuregs[9] [6]), .S0 (n_3040), .Y
       (n_3404));
  MX2X1 g178024(.A (n_386), .B (\cpuregs[9] [7]), .S0 (n_3040), .Y
       (n_3403));
  MX2X1 g178025(.A (n_372), .B (\cpuregs[9] [9]), .S0 (n_3040), .Y
       (n_3402));
  MX2X1 g178026(.A (n_408), .B (\cpuregs[9] [10]), .S0 (n_3040), .Y
       (n_3401));
  MX2X1 g178027(.A (n_418), .B (\cpuregs[9] [8]), .S0 (n_3040), .Y
       (n_3400));
  MX2X1 g178028(.A (n_402), .B (\cpuregs[9] [11]), .S0 (n_3040), .Y
       (n_3399));
  MX2X1 g178029(.A (n_384), .B (\cpuregs[9] [12]), .S0 (n_3040), .Y
       (n_3398));
  MX2X1 g178030(.A (n_388), .B (\cpuregs[9] [13]), .S0 (n_3040), .Y
       (n_3397));
  OAI221X1 g178032(.A0 (n_832), .A1 (n_2943), .B0 (n_2165), .B1
       (n_544), .C0 (n_324), .Y (n_3396));
  AOI22X1 g178033(.A0 (n_2470), .A1 (n_35), .B0 (n_446), .B1 (n_978),
       .Y (n_3469));
  NAND2X1 g178034(.A (n_31), .B (n_1619), .Y (n_3467));
  NAND2X1 g178071(.A (n_2584), .B (n_3175), .Y (n_3466));
  NAND2X1 g178102(.A (n_308), .B (n_3236), .Y (n_3465));
  AND2X2 g178104(.A (n_957), .B (n_3240), .Y (n_333));
  AND2X2 g178105(.A (n_960), .B (n_3244), .Y (n_291));
  AND2X2 g178106(.A (n_964), .B (n_3240), .Y (n_425));
  AND2X2 g178107(.A (n_957), .B (n_3244), .Y (n_424));
  AND2X2 g178108(.A (n_846), .B (n_3240), .Y (n_423));
  AND2X2 g178109(.A (n_957), .B (n_3238), .Y (n_450));
  AND2X2 g178110(.A (n_960), .B (n_3238), .Y (n_462));
  AND2X2 g178111(.A (n_957), .B (n_3237), .Y (n_488));
  AND2X2 g178112(.A (n_964), .B (n_3237), .Y (n_478));
  AND2X2 g178113(.A (n_846), .B (n_3237), .Y (n_486));
  AND2X2 g178114(.A (n_960), .B (n_3237), .Y (n_468));
  AND2X2 g178115(.A (n_964), .B (n_3239), .Y (n_466));
  AND2X2 g178116(.A (n_960), .B (n_3241), .Y (n_464));
  AND2X2 g178117(.A (n_960), .B (n_3242), .Y (n_476));
  AND2X2 g178118(.A (n_846), .B (n_3239), .Y (n_470));
  AND2X2 g178119(.A (n_957), .B (n_3239), .Y (n_484));
  AND2X2 g178120(.A (n_846), .B (n_3241), .Y (n_502));
  AND2X2 g178121(.A (n_957), .B (n_3241), .Y (n_482));
  AND2X2 g178122(.A (n_957), .B (n_3242), .Y (n_500));
  AND2X2 g178123(.A (n_846), .B (n_3242), .Y (n_498));
  AND2X2 g178124(.A (n_960), .B (n_3243), .Y (n_458));
  AND2X2 g178125(.A (n_957), .B (n_3243), .Y (n_480));
  AND2X2 g178126(.A (n_846), .B (n_3243), .Y (n_496));
  AND2X2 g178127(.A (n_964), .B (n_3243), .Y (n_494));
  AND2X2 g178128(.A (n_846), .B (n_3238), .Y (n_448));
  AND2X2 g178129(.A (n_964), .B (n_3241), .Y (n_492));
  AND2X2 g178130(.A (n_964), .B (n_3242), .Y (n_490));
  AND2X2 g178131(.A (n_964), .B (n_3238), .Y (n_452));
  AND2X2 g178132(.A (n_960), .B (n_3239), .Y (n_454));
  AND2X2 g178133(.A (n_960), .B (n_3240), .Y (n_474));
  AND2X2 g178134(.A (n_846), .B (n_3244), .Y (n_456));
  NAND4XL g178135(.A (n_2646), .B (n_2645), .C (n_3013), .D (n_3056),
       .Y (n_3395));
  MX2X1 g178136(.A (n_392), .B (\cpuregs[9] [29]), .S0 (n_3040), .Y
       (n_3394));
  MX2X1 g178137(.A (n_406), .B (\cpuregs[9] [27]), .S0 (n_3040), .Y
       (n_3393));
  MX2X1 g178138(.A (n_370), .B (\cpuregs[9] [30]), .S0 (n_3040), .Y
       (n_3392));
  MX2X1 g178139(.A (n_404), .B (\cpuregs[9] [31]), .S0 (n_3040), .Y
       (n_3391));
  MX2X1 g178140(.A (\cpuregs[17] [1]), .B (n_398), .S0 (n_514), .Y
       (n_3390));
  MX2X1 g178141(.A (\cpuregs[17] [2]), .B (n_366), .S0 (n_514), .Y
       (n_3389));
  MX2X1 g178142(.A (\cpuregs[17] [3]), .B (n_368), .S0 (n_514), .Y
       (n_3388));
  MX2X1 g178143(.A (\cpuregs[17] [4]), .B (n_416), .S0 (n_514), .Y
       (n_3387));
  MX2X1 g178144(.A (\cpuregs[17] [5]), .B (n_394), .S0 (n_514), .Y
       (n_3386));
  MX2X1 g178145(.A (\cpuregs[17] [6]), .B (n_362), .S0 (n_514), .Y
       (n_3385));
  MX2X1 g178146(.A (\cpuregs[17] [7]), .B (n_386), .S0 (n_514), .Y
       (n_3384));
  MX2X1 g178147(.A (\cpuregs[17] [8]), .B (n_418), .S0 (n_514), .Y
       (n_3383));
  MX2X1 g178148(.A (\cpuregs[17] [9]), .B (n_372), .S0 (n_514), .Y
       (n_3382));
  MX2X1 g178149(.A (\cpuregs[17] [10]), .B (n_408), .S0 (n_514), .Y
       (n_3381));
  MX2X1 g178150(.A (\cpuregs[17] [11]), .B (n_402), .S0 (n_514), .Y
       (n_3380));
  MX2X1 g178151(.A (\cpuregs[17] [12]), .B (n_384), .S0 (n_514), .Y
       (n_3379));
  MX2X1 g178152(.A (\cpuregs[17] [13]), .B (n_388), .S0 (n_514), .Y
       (n_3378));
  MX2X1 g178153(.A (\cpuregs[17] [14]), .B (n_374), .S0 (n_514), .Y
       (n_3377));
  MX2X1 g178154(.A (\cpuregs[17] [15]), .B (n_414), .S0 (n_514), .Y
       (n_3376));
  MX2X1 g178155(.A (\cpuregs[17] [16]), .B (n_396), .S0 (n_514), .Y
       (n_3375));
  MX2X1 g178156(.A (\cpuregs[17] [17]), .B (n_412), .S0 (n_514), .Y
       (n_3374));
  MX2X1 g178157(.A (\cpuregs[17] [18]), .B (n_382), .S0 (n_514), .Y
       (n_3373));
  MX2X1 g178158(.A (\cpuregs[17] [20]), .B (n_364), .S0 (n_514), .Y
       (n_3372));
  MX2X1 g178159(.A (\cpuregs[17] [19]), .B (n_1518), .S0 (n_514), .Y
       (n_3371));
  MX2X1 g178160(.A (\cpuregs[17] [21]), .B (n_1515), .S0 (n_514), .Y
       (n_3370));
  MX2X1 g178161(.A (\cpuregs[17] [22]), .B (n_1513), .S0 (n_514), .Y
       (n_3369));
  MX2X1 g178162(.A (\cpuregs[17] [24]), .B (n_378), .S0 (n_514), .Y
       (n_3368));
  MX2X1 g178163(.A (\cpuregs[17] [23]), .B (n_380), .S0 (n_514), .Y
       (n_3367));
  MX2X1 g178164(.A (\cpuregs[17] [25]), .B (n_376), .S0 (n_514), .Y
       (n_3366));
  MX2X1 g178165(.A (\cpuregs[17] [26]), .B (n_400), .S0 (n_514), .Y
       (n_3365));
  MX2X1 g178166(.A (\cpuregs[17] [27]), .B (n_406), .S0 (n_514), .Y
       (n_3364));
  MX2X1 g178167(.A (\cpuregs[17] [28]), .B (n_390), .S0 (n_514), .Y
       (n_3363));
  MX2X1 g178168(.A (\cpuregs[17] [29]), .B (n_392), .S0 (n_514), .Y
       (n_3362));
  MX2X1 g178169(.A (\cpuregs[17] [30]), .B (n_370), .S0 (n_514), .Y
       (n_3361));
  MX2X1 g178170(.A (\cpuregs[17] [31]), .B (n_404), .S0 (n_514), .Y
       (n_3360));
  AOI32X1 g178171(.A0 (n_2997), .A1 (n_2996), .A2 (n_1588), .B0
       (instr_lui), .B1 (n_953), .Y (n_3359));
  MX2X1 g178172(.A (\cpuregs[25] [29]), .B (n_392), .S0 (n_520), .Y
       (n_3358));
  MX2X1 g178173(.A (\cpuregs[25] [25]), .B (n_376), .S0 (n_520), .Y
       (n_3357));
  MX2X1 g178174(.A (\cpuregs[25] [21]), .B (n_1515), .S0 (n_520), .Y
       (n_3356));
  MX2X1 g178175(.A (\cpuregs[25] [1]), .B (n_398), .S0 (n_520), .Y
       (n_3355));
  MX2X1 g178176(.A (\cpuregs[25] [2]), .B (n_366), .S0 (n_520), .Y
       (n_3354));
  MX2X1 g178177(.A (\cpuregs[25] [3]), .B (n_368), .S0 (n_520), .Y
       (n_3353));
  MX2X1 g178178(.A (\cpuregs[25] [4]), .B (n_416), .S0 (n_520), .Y
       (n_3352));
  MX2X1 g178179(.A (\cpuregs[25] [5]), .B (n_394), .S0 (n_520), .Y
       (n_3351));
  MX2X1 g178180(.A (\cpuregs[25] [13]), .B (n_388), .S0 (n_520), .Y
       (n_3350));
  MX2X1 g178181(.A (\cpuregs[25] [6]), .B (n_362), .S0 (n_520), .Y
       (n_3349));
  MX2X1 g178182(.A (\cpuregs[25] [7]), .B (n_386), .S0 (n_520), .Y
       (n_3348));
  MX2X1 g178183(.A (\cpuregs[25] [8]), .B (n_418), .S0 (n_520), .Y
       (n_3347));
  MX2X1 g178184(.A (\cpuregs[25] [9]), .B (n_372), .S0 (n_520), .Y
       (n_3346));
  MX2X1 g178185(.A (\cpuregs[25] [10]), .B (n_408), .S0 (n_520), .Y
       (n_3345));
  MX2X1 g178186(.A (\cpuregs[25] [11]), .B (n_402), .S0 (n_520), .Y
       (n_3344));
  MX2X1 g178187(.A (\cpuregs[25] [12]), .B (n_384), .S0 (n_520), .Y
       (n_3343));
  MX2X1 g178188(.A (\cpuregs[25] [14]), .B (n_374), .S0 (n_520), .Y
       (n_3342));
  MX2X1 g178189(.A (\cpuregs[25] [15]), .B (n_414), .S0 (n_520), .Y
       (n_3341));
  MX2X1 g178190(.A (\cpuregs[25] [16]), .B (n_396), .S0 (n_520), .Y
       (n_3340));
  MX2X1 g178191(.A (\cpuregs[25] [17]), .B (n_412), .S0 (n_520), .Y
       (n_3339));
  MX2X1 g178192(.A (\cpuregs[25] [18]), .B (n_382), .S0 (n_520), .Y
       (n_3338));
  MX2X1 g178193(.A (\cpuregs[25] [19]), .B (n_1518), .S0 (n_520), .Y
       (n_3337));
  MX2X1 g178194(.A (\cpuregs[25] [20]), .B (n_364), .S0 (n_520), .Y
       (n_3336));
  MX2X1 g178195(.A (\cpuregs[25] [22]), .B (n_1513), .S0 (n_520), .Y
       (n_3335));
  MX2X1 g178196(.A (\cpuregs[25] [23]), .B (n_380), .S0 (n_520), .Y
       (n_3334));
  MX2X1 g178197(.A (\cpuregs[25] [24]), .B (n_378), .S0 (n_520), .Y
       (n_3333));
  MX2X1 g178198(.A (\cpuregs[25] [26]), .B (n_400), .S0 (n_520), .Y
       (n_3332));
  MX2X1 g178199(.A (\cpuregs[25] [27]), .B (n_406), .S0 (n_520), .Y
       (n_3331));
  MX2X1 g178200(.A (\cpuregs[25] [28]), .B (n_390), .S0 (n_520), .Y
       (n_3330));
  MX2X1 g178201(.A (\cpuregs[25] [30]), .B (n_370), .S0 (n_520), .Y
       (n_3329));
  MX2X1 g178202(.A (\cpuregs[25] [31]), .B (n_404), .S0 (n_520), .Y
       (n_3328));
  MX2X1 g178203(.A (n_358), .B (\cpuregs[9] [0]), .S0 (n_3040), .Y
       (n_3327));
  MX2X1 g178204(.A (\cpuregs[16] [1]), .B (n_398), .S0 (n_516), .Y
       (n_3326));
  MX2X1 g178205(.A (\cpuregs[16] [2]), .B (n_366), .S0 (n_516), .Y
       (n_3325));
  MX2X1 g178206(.A (\cpuregs[16] [3]), .B (n_368), .S0 (n_516), .Y
       (n_3324));
  MX2X1 g178207(.A (\cpuregs[16] [4]), .B (n_416), .S0 (n_516), .Y
       (n_3323));
  MX2X1 g178208(.A (\cpuregs[16] [5]), .B (n_394), .S0 (n_516), .Y
       (n_3322));
  MX2X1 g178209(.A (\cpuregs[16] [6]), .B (n_362), .S0 (n_516), .Y
       (n_3321));
  MX2X1 g178210(.A (\cpuregs[16] [7]), .B (n_386), .S0 (n_516), .Y
       (n_3320));
  MX2X1 g178211(.A (\cpuregs[16] [8]), .B (n_418), .S0 (n_516), .Y
       (n_3319));
  MX2X1 g178212(.A (\cpuregs[16] [9]), .B (n_372), .S0 (n_516), .Y
       (n_3318));
  MX2X1 g178213(.A (\cpuregs[16] [10]), .B (n_408), .S0 (n_516), .Y
       (n_3317));
  MX2X1 g178214(.A (\cpuregs[16] [11]), .B (n_402), .S0 (n_516), .Y
       (n_3316));
  MX2X1 g178215(.A (\cpuregs[16] [12]), .B (n_384), .S0 (n_516), .Y
       (n_3315));
  MX2X1 g178216(.A (\cpuregs[16] [13]), .B (n_388), .S0 (n_516), .Y
       (n_3314));
  MX2X1 g178217(.A (\cpuregs[16] [14]), .B (n_374), .S0 (n_516), .Y
       (n_3313));
  MX2X1 g178218(.A (\cpuregs[16] [15]), .B (n_414), .S0 (n_516), .Y
       (n_3312));
  MX2X1 g178219(.A (\cpuregs[16] [16]), .B (n_396), .S0 (n_516), .Y
       (n_3311));
  MX2X1 g178220(.A (\cpuregs[16] [17]), .B (n_412), .S0 (n_516), .Y
       (n_3310));
  MX2X1 g178221(.A (\cpuregs[16] [18]), .B (n_382), .S0 (n_516), .Y
       (n_3309));
  MX2X1 g178222(.A (\cpuregs[16] [20]), .B (n_364), .S0 (n_516), .Y
       (n_3308));
  MX2X1 g178223(.A (\cpuregs[16] [19]), .B (n_1518), .S0 (n_516), .Y
       (n_3307));
  MX2X1 g178224(.A (\cpuregs[16] [21]), .B (n_1515), .S0 (n_516), .Y
       (n_3306));
  MX2X1 g178225(.A (\cpuregs[16] [22]), .B (n_1513), .S0 (n_516), .Y
       (n_3305));
  MX2X1 g178226(.A (\cpuregs[16] [23]), .B (n_380), .S0 (n_516), .Y
       (n_3304));
  MX2X1 g178227(.A (\cpuregs[16] [24]), .B (n_378), .S0 (n_516), .Y
       (n_3303));
  MX2X1 g178228(.A (\cpuregs[16] [26]), .B (n_400), .S0 (n_516), .Y
       (n_3302));
  MX2X1 g178229(.A (\cpuregs[16] [27]), .B (n_406), .S0 (n_516), .Y
       (n_3301));
  MX2X1 g178230(.A (\cpuregs[16] [25]), .B (n_376), .S0 (n_516), .Y
       (n_3300));
  MX2X1 g178231(.A (\cpuregs[16] [28]), .B (n_390), .S0 (n_516), .Y
       (n_3299));
  MX2X1 g178232(.A (\cpuregs[16] [29]), .B (n_392), .S0 (n_516), .Y
       (n_3298));
  MX2X1 g178233(.A (\cpuregs[16] [30]), .B (n_370), .S0 (n_516), .Y
       (n_3297));
  MX2X1 g178234(.A (\cpuregs[16] [31]), .B (n_404), .S0 (n_516), .Y
       (n_3296));
  MX2X1 g178235(.A (\cpuregs[24] [1]), .B (n_398), .S0 (n_522), .Y
       (n_3295));
  MX2X1 g178236(.A (\cpuregs[24] [2]), .B (n_366), .S0 (n_522), .Y
       (n_3294));
  MX2X1 g178237(.A (\cpuregs[24] [3]), .B (n_368), .S0 (n_522), .Y
       (n_3293));
  MX2X1 g178238(.A (\cpuregs[24] [4]), .B (n_416), .S0 (n_522), .Y
       (n_3292));
  MX2X1 g178239(.A (\cpuregs[24] [5]), .B (n_394), .S0 (n_522), .Y
       (n_3291));
  MX2X1 g178240(.A (\cpuregs[24] [6]), .B (n_362), .S0 (n_522), .Y
       (n_3290));
  MX2X1 g178241(.A (\cpuregs[24] [7]), .B (n_386), .S0 (n_522), .Y
       (n_3289));
  MX2X1 g178242(.A (\cpuregs[24] [8]), .B (n_418), .S0 (n_522), .Y
       (n_3288));
  MX2X1 g178243(.A (\cpuregs[24] [9]), .B (n_372), .S0 (n_522), .Y
       (n_3287));
  MX2X1 g178244(.A (\cpuregs[24] [10]), .B (n_408), .S0 (n_522), .Y
       (n_3286));
  MX2X1 g178245(.A (\cpuregs[24] [11]), .B (n_402), .S0 (n_522), .Y
       (n_3285));
  MX2X1 g178246(.A (\cpuregs[24] [12]), .B (n_384), .S0 (n_522), .Y
       (n_3284));
  MX2X1 g178247(.A (\cpuregs[24] [13]), .B (n_388), .S0 (n_522), .Y
       (n_3283));
  MX2X1 g178248(.A (\cpuregs[24] [14]), .B (n_374), .S0 (n_522), .Y
       (n_3282));
  MX2X1 g178249(.A (\cpuregs[24] [15]), .B (n_414), .S0 (n_522), .Y
       (n_3281));
  MX2X1 g178250(.A (\cpuregs[24] [16]), .B (n_396), .S0 (n_522), .Y
       (n_3280));
  MX2X1 g178251(.A (\cpuregs[24] [17]), .B (n_412), .S0 (n_522), .Y
       (n_3279));
  MX2X1 g178252(.A (\cpuregs[24] [18]), .B (n_382), .S0 (n_522), .Y
       (n_3278));
  MX2X1 g178253(.A (\cpuregs[24] [19]), .B (n_1518), .S0 (n_522), .Y
       (n_3277));
  MX2X1 g178254(.A (\cpuregs[24] [20]), .B (n_364), .S0 (n_522), .Y
       (n_3276));
  MX2X1 g178255(.A (\cpuregs[24] [22]), .B (n_1513), .S0 (n_522), .Y
       (n_3275));
  MX2X1 g178256(.A (\cpuregs[24] [23]), .B (n_380), .S0 (n_522), .Y
       (n_3274));
  MX2X1 g178257(.A (\cpuregs[24] [24]), .B (n_378), .S0 (n_522), .Y
       (n_3273));
  MX2X1 g178258(.A (\cpuregs[24] [25]), .B (n_376), .S0 (n_522), .Y
       (n_3272));
  MX2X1 g178259(.A (\cpuregs[24] [26]), .B (n_400), .S0 (n_522), .Y
       (n_3271));
  MX2X1 g178260(.A (\cpuregs[24] [27]), .B (n_406), .S0 (n_522), .Y
       (n_3270));
  MX2X1 g178261(.A (\cpuregs[24] [28]), .B (n_390), .S0 (n_522), .Y
       (n_3269));
  MX2X1 g178262(.A (\cpuregs[24] [29]), .B (n_392), .S0 (n_522), .Y
       (n_3268));
  MX2X1 g178263(.A (\cpuregs[24] [30]), .B (n_370), .S0 (n_522), .Y
       (n_3267));
  MX2X1 g178264(.A (\cpuregs[24] [31]), .B (n_404), .S0 (n_522), .Y
       (n_3266));
  MX2X1 g178265(.A (\cpuregs[24] [21]), .B (n_1515), .S0 (n_522), .Y
       (n_3265));
  MX2X1 g178266(.A (\cpuregs[17] [0]), .B (n_358), .S0 (n_514), .Y
       (n_3264));
  MX2X1 g178267(.A (\cpuregs[25] [0]), .B (n_358), .S0 (n_520), .Y
       (n_3263));
  MX2X1 g178268(.A (\cpuregs[16] [0]), .B (n_358), .S0 (n_516), .Y
       (n_3262));
  MX2X1 g178269(.A (\cpuregs[24] [0]), .B (n_358), .S0 (n_522), .Y
       (n_3261));
  MX2X1 g178270(.A (mem_rdata_q[10]), .B (n_503), .S0 (n_35), .Y
       (n_3260));
  MX2X1 g178271(.A (mem_rdata_q[11]), .B (n_440), .S0 (n_35), .Y
       (n_3259));
  OAI22X1 g178272(.A0 (n_679), .A1 (n_3070), .B0 (n_683), .B1 (n_2422),
       .Y (n_3258));
  AOI32X1 g178273(.A0 (n_2144), .A1 (n_2604), .A2 (n_35), .B0 (n_334),
       .B1 (n_2436), .Y (n_3257));
  NAND4XL g178274(.A (n_2881), .B (n_2856), .C (n_3011), .D (n_3048),
       .Y (n_3256));
  NAND4XL g178275(.A (n_2710), .B (n_2709), .C (n_3010), .D (n_3055),
       .Y (n_3255));
  MX2X1 g178276(.A (n_390), .B (\cpuregs[9] [28]), .S0 (n_3040), .Y
       (n_3254));
  INVX1 g178277(.A (n_3252), .Y (n_3253));
  INVX1 g178278(.A (n_3247), .Y (n_3248));
  INVX1 g178279(.A (n_3245), .Y (n_3246));
  MX2X1 g178281(.A (\cpuregs[1] [2]), .B (n_366), .S0 (n_508), .Y
       (n_3210));
  MX2X1 g178282(.A (\cpuregs[1] [1]), .B (n_398), .S0 (n_508), .Y
       (n_3209));
  MX2X1 g178283(.A (\cpuregs[8] [31]), .B (n_404), .S0 (n_506), .Y
       (n_3208));
  MX2X1 g178284(.A (\cpuregs[8] [30]), .B (n_370), .S0 (n_506), .Y
       (n_3207));
  MX2X1 g178285(.A (\cpuregs[8] [29]), .B (n_392), .S0 (n_506), .Y
       (n_3206));
  MX2X1 g178286(.A (\cpuregs[8] [28]), .B (n_390), .S0 (n_506), .Y
       (n_3205));
  MX2X1 g178287(.A (\cpuregs[8] [27]), .B (n_406), .S0 (n_506), .Y
       (n_3204));
  MX2X1 g178288(.A (\cpuregs[8] [26]), .B (n_400), .S0 (n_506), .Y
       (n_3203));
  MX2X1 g178289(.A (\cpuregs[8] [25]), .B (n_376), .S0 (n_506), .Y
       (n_3202));
  MX2X1 g178290(.A (\cpuregs[8] [24]), .B (n_378), .S0 (n_506), .Y
       (n_3201));
  MX2X1 g178291(.A (\cpuregs[8] [21]), .B (n_1515), .S0 (n_506), .Y
       (n_3200));
  MX2X1 g178292(.A (\cpuregs[8] [23]), .B (n_380), .S0 (n_506), .Y
       (n_3199));
  MX2X1 g178293(.A (\cpuregs[8] [22]), .B (n_1513), .S0 (n_506), .Y
       (n_3198));
  MX2X1 g178294(.A (\cpuregs[8] [20]), .B (n_364), .S0 (n_506), .Y
       (n_3197));
  MX2X1 g178295(.A (\cpuregs[8] [19]), .B (n_1518), .S0 (n_506), .Y
       (n_3196));
  MX2X1 g178296(.A (\cpuregs[8] [18]), .B (n_382), .S0 (n_506), .Y
       (n_3195));
  MX2X1 g178297(.A (\cpuregs[8] [17]), .B (n_412), .S0 (n_506), .Y
       (n_3194));
  NOR2X1 g178298(.A (n_2347), .B (n_3019), .Y (n_3193));
  MX2X1 g178299(.A (\cpuregs[8] [15]), .B (n_414), .S0 (n_506), .Y
       (n_3192));
  MX2X1 g178300(.A (\cpuregs[8] [16]), .B (n_396), .S0 (n_506), .Y
       (n_3191));
  MX2X1 g178301(.A (\cpuregs[8] [14]), .B (n_374), .S0 (n_506), .Y
       (n_3190));
  MX2X1 g178302(.A (\cpuregs[8] [13]), .B (n_388), .S0 (n_506), .Y
       (n_3189));
  MX2X1 g178303(.A (\cpuregs[8] [12]), .B (n_384), .S0 (n_506), .Y
       (n_3188));
  MX2X1 g178304(.A (\cpuregs[8] [11]), .B (n_402), .S0 (n_506), .Y
       (n_3187));
  MX2X1 g178305(.A (\cpuregs[8] [9]), .B (n_372), .S0 (n_506), .Y
       (n_3186));
  MX2X1 g178306(.A (\cpuregs[8] [10]), .B (n_408), .S0 (n_506), .Y
       (n_3185));
  MX2X1 g178307(.A (\cpuregs[8] [2]), .B (n_366), .S0 (n_506), .Y
       (n_3184));
  MX2X1 g178308(.A (\cpuregs[8] [7]), .B (n_386), .S0 (n_506), .Y
       (n_3183));
  MX2X1 g178309(.A (\cpuregs[8] [6]), .B (n_362), .S0 (n_506), .Y
       (n_3182));
  MX2X1 g178310(.A (\cpuregs[8] [5]), .B (n_394), .S0 (n_506), .Y
       (n_3181));
  MX2X1 g178311(.A (\cpuregs[8] [4]), .B (n_416), .S0 (n_506), .Y
       (n_3180));
  MX2X1 g178312(.A (\cpuregs[8] [3]), .B (n_368), .S0 (n_506), .Y
       (n_3179));
  MX2X1 g178313(.A (\cpuregs[8] [1]), .B (n_398), .S0 (n_506), .Y
       (n_3178));
  MX2X1 g178314(.A (\cpuregs[8] [8]), .B (n_418), .S0 (n_506), .Y
       (n_3177));
  OAI211X1 g178315(.A0 (n_603), .A1 (n_2326), .B0 (n_542), .C0 (n_314),
       .Y (n_3176));
  AOI221X1 g178316(.A0 (n_317), .A1 (n_13), .B0 (n_2439), .B1 (n_1588),
       .C0 (n_3046), .Y (n_3175));
  NOR2X1 g178317(.A (n_17), .B (n_3066), .Y (n_3174));
  OAI31X1 g178318(.A0 (n_317), .A1 (n_2320), .A2 (n_2600), .B0
       (n_2534), .Y (n_3173));
  OAI211X1 g178319(.A0 (n_764), .A1 (n_2326), .B0 (n_1628), .C0
       (n_314), .Y (n_3172));
  NAND4XL g178320(.A (n_635), .B (n_714), .C
       (\genblk2.pcpi_div_minus_2470_59_n_502 ), .D (n_2571), .Y
       (n_3171));
  AOI221X1 g178321(.A0 (n_334), .A1 (n_2608), .B0 (is_alu_reg_reg), .B1
       (n_953), .C0 (n_3009), .Y (n_3170));
  NAND4XL g178322(.A (n_1196), .B (n_1195), .C (n_1352), .D (n_2567),
       .Y (n_3169));
  AOI22X1 g178323(.A0 (n_852), .A1 (n_2611), .B0 (n_1731), .B1
       (n_1184), .Y (n_3168));
  AOI211XL g178324(.A0 (\cpuregs[18] [1]), .A1 (n_10), .B0 (n_2353),
       .C0 (n_2948), .Y (n_3167));
  AOI211XL g178325(.A0 (\cpuregs[28] [0]), .A1 (n_9), .B0 (n_2352), .C0
       (n_2949), .Y (n_3166));
  OAI2BB1X1 g178326(.A0N (n_2822), .A1N (n_1619), .B0 (n_2605), .Y
       (n_3252));
  NOR4X1 g178327(.A (mem_rdata_q[24]), .B (mem_rdata_q[15]), .C
       (n_586), .D (n_2597), .Y (n_3251));
  NAND3X1 g178329(.A (n_18), .B (n_2996), .C (n_1588), .Y (n_3250));
  NOR2X1 g178331(.A (n_3066), .B (n_2436), .Y (n_3249));
  NAND4BX1 g178332(.AN (n_3020), .B (n_2034), .C (n_2033), .D (n_2555),
       .Y (n_3247));
  NAND4BX1 g178333(.AN (n_3021), .B (n_2064), .C (n_2026), .D (n_2558),
       .Y (n_3245));
  NOR2X1 g178334(.A (decoded_rs1[4]), .B (n_3072), .Y (n_3244));
  AND2X1 g178336(.A (n_3074), .B (decoded_rs1[4]), .Y (n_3243));
  NOR2X1 g178337(.A (n_574), .B (n_20), .Y (n_3242));
  NOR2X1 g178338(.A (n_574), .B (n_3073), .Y (n_3241));
  NOR2X1 g178339(.A (decoded_rs1[4]), .B (n_3073), .Y (n_3240));
  AND2X1 g178340(.A (n_3074), .B (n_574), .Y (n_3239));
  NOR2X1 g178341(.A (decoded_rs1[4]), .B (n_20), .Y (n_3238));
  NOR2X1 g178342(.A (n_574), .B (n_3072), .Y (n_3237));
  NAND2X1 g178345(.A (n_445), .B (n_308), .Y (n_3236));
  NAND2X1 g178346(.A (n_317), .B (n_696), .Y (n_329));
  AND2X2 g178348(.A (n_847), .B (n_3041), .Y (n_536));
  OR2X2 g178349(.A (n_848), .B (n_347), .Y (n_3233));
  AND2X2 g178350(.A (n_965), .B (n_19), .Y (n_510));
  AND2X2 g178351(.A (n_847), .B (n_19), .Y (n_512));
  AND2X2 g178352(.A (n_845), .B (n_19), .Y (n_518));
  OR2X2 g178353(.A (n_848), .B (n_21), .Y (n_3229));
  AND2X2 g178354(.A (n_290), .B (n_19), .Y (n_528));
  AND2X2 g178355(.A (n_290), .B (n_3041), .Y (n_534));
  OR2X2 g178356(.A (n_671), .B (n_21), .Y (n_3226));
  OR2X2 g178357(.A (n_848), .B (n_3068), .Y (n_3225));
  AND2X2 g178358(.A (n_290), .B (n_3067), .Y (n_526));
  AND2X2 g178359(.A (n_290), .B (n_695), .Y (n_524));
  AND2X2 g178360(.A (n_845), .B (n_3041), .Y (n_532));
  OR2X2 g178361(.A (n_966), .B (n_347), .Y (n_3221));
  OR2X2 g178362(.A (n_671), .B (n_3069), .Y (n_3220));
  OR2X2 g178363(.A (n_966), .B (n_3069), .Y (n_3219));
  OR2X2 g178364(.A (n_966), .B (n_21), .Y (n_3218));
  OR2X2 g178365(.A (n_844), .B (n_21), .Y (n_3217));
  OR2X2 g178366(.A (n_844), .B (n_3069), .Y (n_3216));
  OR2X2 g178367(.A (n_966), .B (n_3068), .Y (n_3215));
  OR2X2 g178368(.A (n_844), .B (n_347), .Y (n_3214));
  OR2X2 g178369(.A (n_844), .B (n_3068), .Y (n_3213));
  OR2X2 g178370(.A (n_848), .B (n_3069), .Y (n_3212));
  AND2X2 g178371(.A (n_965), .B (n_3041), .Y (n_530));
  NAND4XL g178373(.A (n_2831), .B (n_2901), .C (n_2833), .D (n_2832),
       .Y (n_3165));
  MX2X1 g178374(.A (\cpuregs[1] [4]), .B (n_416), .S0 (n_508), .Y
       (n_3164));
  MX2X1 g178375(.A (\cpuregs[1] [5]), .B (n_394), .S0 (n_508), .Y
       (n_3163));
  MX2X1 g178376(.A (\cpuregs[1] [6]), .B (n_362), .S0 (n_508), .Y
       (n_3162));
  MX2X1 g178377(.A (\cpuregs[1] [7]), .B (n_386), .S0 (n_508), .Y
       (n_3161));
  MX2X1 g178378(.A (\cpuregs[1] [8]), .B (n_418), .S0 (n_508), .Y
       (n_3160));
  MX2X1 g178379(.A (\cpuregs[1] [9]), .B (n_372), .S0 (n_508), .Y
       (n_3159));
  MX2X1 g178380(.A (\cpuregs[1] [10]), .B (n_408), .S0 (n_508), .Y
       (n_3158));
  MX2X1 g178381(.A (\cpuregs[1] [11]), .B (n_402), .S0 (n_508), .Y
       (n_3157));
  MX2X1 g178382(.A (\cpuregs[1] [13]), .B (n_388), .S0 (n_508), .Y
       (n_3156));
  MX2X1 g178383(.A (\cpuregs[1] [14]), .B (n_374), .S0 (n_508), .Y
       (n_3155));
  MX2X1 g178384(.A (\cpuregs[1] [15]), .B (n_414), .S0 (n_508), .Y
       (n_3154));
  MX2X1 g178385(.A (\cpuregs[1] [12]), .B (n_384), .S0 (n_508), .Y
       (n_3153));
  MX2X1 g178386(.A (\cpuregs[1] [16]), .B (n_396), .S0 (n_508), .Y
       (n_3152));
  MX2X1 g178387(.A (\cpuregs[1] [17]), .B (n_412), .S0 (n_508), .Y
       (n_3151));
  MX2X1 g178388(.A (\cpuregs[1] [18]), .B (n_382), .S0 (n_508), .Y
       (n_3150));
  MX2X1 g178389(.A (\cpuregs[1] [19]), .B (n_1518), .S0 (n_508), .Y
       (n_3149));
  MX2X1 g178390(.A (\cpuregs[1] [20]), .B (n_364), .S0 (n_508), .Y
       (n_3148));
  MX2X1 g178391(.A (\cpuregs[1] [21]), .B (n_1515), .S0 (n_508), .Y
       (n_3147));
  MX2X1 g178392(.A (\cpuregs[1] [22]), .B (n_1513), .S0 (n_508), .Y
       (n_3146));
  MX2X1 g178393(.A (\cpuregs[1] [23]), .B (n_380), .S0 (n_508), .Y
       (n_3145));
  MX2X1 g178394(.A (\cpuregs[1] [25]), .B (n_376), .S0 (n_508), .Y
       (n_3144));
  MX2X1 g178395(.A (\cpuregs[1] [24]), .B (n_378), .S0 (n_508), .Y
       (n_3143));
  MX2X1 g178396(.A (\cpuregs[1] [26]), .B (n_400), .S0 (n_508), .Y
       (n_3142));
  MX2X1 g178397(.A (\cpuregs[1] [27]), .B (n_406), .S0 (n_508), .Y
       (n_3141));
  MX2X1 g178398(.A (\cpuregs[1] [28]), .B (n_390), .S0 (n_508), .Y
       (n_3140));
  MX2X1 g178399(.A (\cpuregs[1] [30]), .B (n_370), .S0 (n_508), .Y
       (n_3139));
  MX2X1 g178400(.A (\cpuregs[1] [31]), .B (n_404), .S0 (n_508), .Y
       (n_3138));
  MX2X1 g178401(.A (\cpuregs[1] [29]), .B (n_392), .S0 (n_508), .Y
       (n_3137));
  MX2X1 g178402(.A (\cpuregs[8] [0]), .B (n_358), .S0 (n_506), .Y
       (n_3136));
  MX2X1 g178403(.A (\cpuregs[1] [0]), .B (n_358), .S0 (n_508), .Y
       (n_3135));
  NAND4XL g178404(.A (n_2811), .B (n_2813), .C (n_2812), .D (n_2814),
       .Y (n_3134));
  NAND4XL g178405(.A (n_2961), .B (n_2960), .C (n_2915), .D (n_2959),
       .Y (n_3133));
  NAND4XL g178406(.A (n_2954), .B (n_2952), .C (n_2953), .D (n_2951),
       .Y (n_3132));
  NAND4XL g178407(.A (n_2648), .B (n_2913), .C (n_2650), .D (n_2649),
       .Y (n_3131));
  NAND4XL g178408(.A (n_2848), .B (n_2910), .C (n_2894), .D (n_2849),
       .Y (n_3130));
  NAND4XL g178409(.A (n_2886), .B (n_2889), .C (n_2888), .D (n_2940),
       .Y (n_3129));
  NAND4XL g178410(.A (n_2883), .B (n_2935), .C (n_2885), .D (n_2884),
       .Y (n_3128));
  NAND4XL g178411(.A (n_2879), .B (n_2882), .C (n_2880), .D (n_2941),
       .Y (n_3127));
  NAND4XL g178412(.A (n_2874), .B (n_2875), .C (n_2617), .D (n_2616),
       .Y (n_3126));
  NAND4XL g178413(.A (n_2868), .B (n_2870), .C (n_2869), .D (n_2985),
       .Y (n_3125));
  NAND4XL g178414(.A (n_2858), .B (n_2861), .C (n_2860), .D (n_2859),
       .Y (n_3124));
  NAND4XL g178415(.A (n_2852), .B (n_2854), .C (n_2853), .D (n_2892),
       .Y (n_3123));
  NAND4XL g178416(.A (n_2845), .B (n_2900), .C (n_2846), .D (n_2895),
       .Y (n_3122));
  NAND4XL g178417(.A (n_2838), .B (n_2840), .C (n_2839), .D (n_2841),
       .Y (n_3121));
  NAND4XL g178418(.A (n_2898), .B (n_2835), .C (n_2834), .D (n_2907),
       .Y (n_3120));
  MX2X1 g178419(.A (\cpuregs[1] [3]), .B (n_368), .S0 (n_508), .Y
       (n_3119));
  NAND4XL g178420(.A (n_2927), .B (n_2830), .C (n_2829), .D (n_2902),
       .Y (n_3118));
  NAND4XL g178421(.A (n_2826), .B (n_2828), .C (n_2827), .D (n_2905),
       .Y (n_3117));
  NAND4XL g178422(.A (n_2893), .B (n_2823), .C (n_2909), .D (n_2908),
       .Y (n_3116));
  NAND4XL g178423(.A (n_2971), .B (n_2963), .C (n_2965), .D (n_2918),
       .Y (n_3115));
  NAND4XL g178424(.A (n_2979), .B (n_2977), .C (n_2978), .D (n_2920),
       .Y (n_3114));
  NAND4XL g178425(.A (n_2922), .B (n_2982), .C (n_2983), .D (n_2921),
       .Y (n_3113));
  NAND4XL g178426(.A (n_2988), .B (n_2987), .C (n_2925), .D (n_2986),
       .Y (n_3112));
  NAND4XL g178427(.A (n_2992), .B (n_2990), .C (n_2991), .D (n_2931),
       .Y (n_3111));
  NAND4XL g178428(.A (n_2817), .B (n_2818), .C (n_2934), .D (n_2933),
       .Y (n_3110));
  NAND4XL g178429(.A (n_2808), .B (n_2809), .C (n_2939), .D (n_2938),
       .Y (n_3109));
  NAND4XL g178430(.A (n_2802), .B (n_2804), .C (n_2803), .D (n_2942),
       .Y (n_3108));
  NAND4XL g178431(.A (n_2800), .B (n_2896), .C (n_2638), .D (n_2801),
       .Y (n_3107));
  NAND4XL g178432(.A (n_2871), .B (n_2786), .C (n_2873), .D (n_2872),
       .Y (n_3106));
  NAND4XL g178433(.A (n_2796), .B (n_2799), .C (n_2798), .D (n_2797),
       .Y (n_3105));
  NAND4XL g178434(.A (n_2790), .B (n_2792), .C (n_2791), .D (n_2793),
       .Y (n_3104));
  NAND4XL g178435(.A (n_2782), .B (n_2784), .C (n_2783), .D (n_2785),
       .Y (n_3103));
  NAND4XL g178436(.A (n_2777), .B (n_2779), .C (n_2778), .D (n_2911),
       .Y (n_3102));
  NAND4XL g178437(.A (n_2770), .B (n_2772), .C (n_2771), .D (n_2773),
       .Y (n_3101));
  NAND4XL g178438(.A (n_2764), .B (n_2766), .C (n_2765), .D (n_2767),
       .Y (n_3100));
  NAND4XL g178439(.A (n_2757), .B (n_2760), .C (n_2759), .D (n_2758),
       .Y (n_3099));
  NAND4XL g178440(.A (n_2752), .B (n_2754), .C (n_2753), .D (n_2916),
       .Y (n_3098));
  NAND4XL g178441(.A (n_2745), .B (n_2747), .C (n_2746), .D (n_2748),
       .Y (n_3097));
  NAND4XL g178442(.A (n_2739), .B (n_2741), .C (n_2740), .D (n_2742),
       .Y (n_3096));
  NAND4XL g178443(.A (n_2732), .B (n_2734), .C (n_2733), .D (n_2735),
       .Y (n_3095));
  NAND4XL g178444(.A (n_2726), .B (n_2728), .C (n_2727), .D (n_2929),
       .Y (n_3094));
  NAND4XL g178445(.A (n_2723), .B (n_2630), .C (n_2725), .D (n_2724),
       .Y (n_3093));
  NAND4XL g178446(.A (n_2720), .B (n_2722), .C (n_2721), .D (n_2928),
       .Y (n_3092));
  NAND4XL g178447(.A (n_2712), .B (n_2864), .C (n_2821), .D (n_2713),
       .Y (n_3091));
  NAND4XL g178448(.A (n_2703), .B (n_2705), .C (n_2704), .D (n_2706),
       .Y (n_3090));
  NAND4XL g178449(.A (n_2696), .B (n_2698), .C (n_2697), .D (n_2699),
       .Y (n_3089));
  NAND4XL g178450(.A (n_2690), .B (n_2692), .C (n_2691), .D (n_2865),
       .Y (n_3088));
  NAND4XL g178451(.A (n_2686), .B (n_2689), .C (n_2688), .D (n_2687),
       .Y (n_3087));
  NAND4XL g178452(.A (n_2682), .B (n_2685), .C (n_2684), .D (n_2683),
       .Y (n_3086));
  NAND4XL g178453(.A (n_2677), .B (n_2679), .C (n_2678), .D (n_2899),
       .Y (n_3085));
  NAND4XL g178454(.A (n_2670), .B (n_2672), .C (n_2671), .D (n_2673),
       .Y (n_3084));
  NAND4XL g178455(.A (n_2663), .B (n_2665), .C (n_2664), .D (n_2666),
       .Y (n_3083));
  NAND4XL g178456(.A (n_2659), .B (n_2662), .C (n_2661), .D (n_2660),
       .Y (n_3082));
  NAND4XL g178457(.A (n_2932), .B (n_2658), .C (n_2657), .D (n_2656),
       .Y (n_3081));
  NAND4XL g178458(.A (n_2639), .B (n_2641), .C (n_2640), .D (n_2642),
       .Y (n_3080));
  NAND4XL g178459(.A (n_2631), .B (n_2634), .C (n_2633), .D (n_2632),
       .Y (n_3079));
  NAND4XL g178460(.A (n_2625), .B (n_2627), .C (n_2626), .D (n_2930),
       .Y (n_3078));
  NAND4XL g178461(.A (n_2618), .B (n_2620), .C (n_2619), .D (n_2621),
       .Y (n_3077));
  OAI31X1 g178462(.A0 (mem_rdata_latched[0]), .A1 (n_692), .A2 (n_335),
       .B0 (n_3014), .Y (n_3076));
  AOI222X1 g178463(.A0 (n_429), .A1 (n_673), .B0 (is_lb_lh_lw_lbu_lhu),
       .B1 (n_953), .C0 (n_2440), .C1 (n_419), .Y (n_3075));
  INVX1 g178465(.A (n_3070), .Y (n_3071));
  INVX1 g178466(.A (n_3068), .Y (n_3067));
  INVX1 g178467(.A (n_3066), .Y (n_3065));
  AOI221X1 g178469(.A0 (\cpuregs[1] [16]), .A1 (n_552), .B0
       (\cpuregs[31] [16]), .B1 (n_2499), .C0 (n_1764), .Y (n_3059));
  AOI221X1 g178470(.A0 (\cpuregs[31] [17]), .A1 (n_2499), .B0
       (\reg_op2[17]_9686 ), .B1 (n_832), .C0 (n_2805), .Y (n_3058));
  AOI221X1 g178471(.A0 (\cpuregs[1] [30]), .A1 (n_552), .B0
       (\cpuregs[31] [30]), .B1 (n_2499), .C0 (n_1776), .Y (n_3057));
  AOI221X1 g178472(.A0 (\cpuregs[8] [29]), .A1 (n_2494), .B0
       (\cpuregs[11] [29]), .B1 (n_2497), .C0 (n_2647), .Y (n_3056));
  AOI221X1 g178473(.A0 (\cpuregs[10] [24]), .A1 (n_2520), .B0
       (\cpuregs[13] [24]), .B1 (n_2498), .C0 (n_2711), .Y (n_3055));
  AOI221X1 g178474(.A0 (\cpuregs[31] [23]), .A1 (n_2499), .B0
       (\reg_op2[23]_9692 ), .B1 (n_832), .C0 (n_2729), .Y (n_3054));
  AOI221X1 g178475(.A0 (\cpuregs[1] [22]), .A1 (n_552), .B0
       (\cpuregs[31] [22]), .B1 (n_2499), .C0 (n_1759), .Y (n_3053));
  OR4X1 g178476(.A (\genblk2.pcpi_div_quotient_msk [16]), .B
       (\genblk2.pcpi_div_quotient_msk [15]), .C
       (\genblk2.pcpi_div_quotient_msk [14]), .D (n_2516), .Y (n_3052));
  OAI2BB1X1 g178477(.A0N (n_6535), .A1N (n_2595), .B0 (n_6538), .Y
       (n_3051));
  AOI221X1 g178478(.A0 (\cpuregs[1] [21]), .A1 (n_552), .B0
       (\cpuregs[31] [21]), .B1 (n_2499), .C0 (n_1760), .Y (n_3050));
  AOI221X1 g178479(.A0 (\cpuregs[1] [19]), .A1 (n_552), .B0
       (\cpuregs[31] [19]), .B1 (n_2499), .C0 (n_1762), .Y (n_3049));
  AOI221X1 g178480(.A0 (\cpuregs[8] [7]), .A1 (n_2494), .B0
       (\cpuregs[7] [7]), .B1 (n_12), .C0 (n_2857), .Y (n_3048));
  NOR2X1 g178481(.A (n_544), .B (n_2944), .Y (n_3047));
  NOR2X1 g178484(.A (decoded_rs1[1]), .B (n_3002), .Y (n_3074));
  NAND2X1 g178485(.A (decoded_rs1[1]), .B (n_3003), .Y (n_3073));
  NAND2BX1 g178486(.AN (decoded_rs1[1]), .B (n_3003), .Y (n_3072));
  NOR2X1 g178493(.A (n_17), .B (n_2998), .Y (n_3070));
  NAND2X1 g178498(.A (n_638), .B (n_3001), .Y (n_3069));
  NAND2X1 g178499(.A (latched_rd[2]), .B (n_3004), .Y (n_3068));
  NOR2BX1 g178501(.AN (n_18), .B (n_1590), .Y (n_3066));
  NAND2X1 g178502(.A (n_2997), .B (n_1589), .Y (n_308));
  AND2X2 g178503(.A (n_845), .B (n_2999), .Y (n_516));
  AND2X2 g178504(.A (n_290), .B (n_2999), .Y (n_522));
  AND2X2 g178505(.A (n_290), .B (n_3000), .Y (n_520));
  AND2X2 g178506(.A (n_845), .B (n_3000), .Y (n_514));
  INVX1 g178507(.A (n_3045), .Y (n_3046));
  OAI211X1 g178509(.A0 (n_130), .A1 (n_667), .B0 (n_2563), .C0
       (n_2448), .Y (n_3039));
  AOI221X1 g178510(.A0 (\cpuregs[1] [14]), .A1 (n_552), .B0
       (\cpuregs[31] [14]), .B1 (n_2499), .C0 (n_1775), .Y (n_3038));
  AOI221X1 g178511(.A0 (\cpuregs[1] [9]), .A1 (n_552), .B0
       (\cpuregs[31] [9]), .B1 (n_2499), .C0 (n_1767), .Y (n_3037));
  AOI221X1 g178512(.A0 (\cpuregs[1] [8]), .A1 (n_552), .B0
       (\cpuregs[31] [8]), .B1 (n_2499), .C0 (n_1773), .Y (n_3036));
  AOI221X1 g178513(.A0 (\cpuregs[31] [5]), .A1 (n_2499), .B0
       (\reg_op2[5]_9674 ), .B1 (n_832), .C0 (n_2890), .Y (n_3035));
  AOI221X1 g178514(.A0 (\cpuregs[31] [6]), .A1 (n_2499), .B0
       (\reg_op2[6]_9675 ), .B1 (n_832), .C0 (n_2876), .Y (n_3034));
  AOI221X1 g178515(.A0 (\cpuregs[31] [10]), .A1 (n_2499), .B0
       (\reg_op2[10]_9679 ), .B1 (n_832), .C0 (n_2836), .Y (n_3033));
  AOI221X1 g178516(.A0 (\cpuregs[1] [11]), .A1 (n_552), .B0
       (\cpuregs[31] [11]), .B1 (n_2499), .C0 (n_1766), .Y (n_3032));
  AOI221X1 g178517(.A0 (\cpuregs[1] [12]), .A1 (n_552), .B0
       (\cpuregs[31] [12]), .B1 (n_2499), .C0 (n_1769), .Y (n_3031));
  AOI221X1 g178518(.A0 (\cpuregs[1] [13]), .A1 (n_552), .B0
       (\cpuregs[31] [13]), .B1 (n_2499), .C0 (n_1765), .Y (n_3030));
  AOI221X1 g178519(.A0 (\cpuregs[1] [15]), .A1 (n_552), .B0
       (\cpuregs[31] [15]), .B1 (n_2499), .C0 (n_1778), .Y (n_3029));
  AOI221X1 g178520(.A0 (\cpuregs[1] [18]), .A1 (n_552), .B0
       (\cpuregs[31] [18]), .B1 (n_2499), .C0 (n_1763), .Y (n_3028));
  AOI221X1 g178521(.A0 (\cpuregs[1] [20]), .A1 (n_552), .B0
       (\cpuregs[31] [20]), .B1 (n_2499), .C0 (n_1761), .Y (n_3027));
  AOI221X1 g178522(.A0 (\cpuregs[1] [25]), .A1 (n_552), .B0
       (\cpuregs[31] [25]), .B1 (n_2499), .C0 (n_1758), .Y (n_3026));
  AOI221X1 g178523(.A0 (\cpuregs[31] [26]), .A1 (n_2499), .B0
       (\reg_op2[26]_9695 ), .B1 (n_832), .C0 (n_2693), .Y (n_3025));
  AOI221X1 g178524(.A0 (\cpuregs[1] [27]), .A1 (n_552), .B0
       (\cpuregs[31] [27]), .B1 (n_2499), .C0 (n_1757), .Y (n_3024));
  AOI221X1 g178525(.A0 (\cpuregs[31] [28]), .A1 (n_2499), .B0
       (\reg_op2[28]_9697 ), .B1 (n_832), .C0 (n_2667), .Y (n_3023));
  AOI221X1 g178526(.A0 (\cpuregs[1] [31]), .A1 (n_552), .B0
       (\cpuregs[31] [31]), .B1 (n_2499), .C0 (n_1782), .Y (n_3022));
  NAND4XL g178527(.A (n_2022), .B (n_2023), .C (n_2065), .D (n_2575),
       .Y (n_3021));
  NAND4XL g178528(.A (n_2029), .B (n_2060), .C (n_2061), .D (n_2576),
       .Y (n_3020));
  NAND4XL g178529(.A (n_2013), .B (n_2071), .C (n_2014), .D (n_2574),
       .Y (n_3019));
  OAI32X1 g178530(.A0 (n_622), .A1 (n_537), .A2 (n_2509), .B0 (n_599),
       .B1 (n_538), .Y (n_3018));
  OAI211X1 g178531(.A0 (n_652), .A1 (n_667), .B0 (n_2609), .C0
       (n_2425), .Y (n_3017));
  OAI2BB1X1 g178532(.A0N (instr_auipc), .A1N (n_953), .B0 (n_2614), .Y
       (n_3016));
  AOI22X1 g178533(.A0 (n_2572), .A1 (n_1588), .B0 (n_692), .B1 (n_419),
       .Y (n_3015));
  AOI22X1 g178534(.A0 (n_679), .A1 (n_2608), .B0 (is_sb_sh_sw), .B1
       (n_953), .Y (n_3014));
  AOI222X1 g178535(.A0 (\cpuregs[1] [29]), .A1 (n_552), .B0
       (\cpuregs[14] [29]), .B1 (n_2531), .C0 (\cpuregs[9] [29]), .C1
       (n_2526), .Y (n_3013));
  OAI32X1 g178536(.A0 (n_729), .A1 (n_537), .A2 (n_2509), .B0 (n_767),
       .B1 (n_538), .Y (n_3012));
  AOI222X1 g178537(.A0 (\cpuregs[1] [7]), .A1 (n_552), .B0
       (\cpuregs[14] [7]), .B1 (n_2531), .C0 (\cpuregs[9] [7]), .C1
       (n_2526), .Y (n_3011));
  AOI222X1 g178538(.A0 (\cpuregs[1] [24]), .A1 (n_552), .B0
       (\cpuregs[14] [24]), .B1 (n_2531), .C0 (\cpuregs[7] [24]), .C1
       (n_12), .Y (n_3010));
  NAND3X1 g178539(.A (n_2600), .B (n_2995), .C (n_13), .Y (n_3045));
  NAND3X1 g178541(.A (n_2440), .B (n_2600), .C (n_1619), .Y (n_3044));
  OAI211X1 g178542(.A0 (n_11741), .A1 (n_2532), .B0 (n_2605), .C0
       (n_2602), .Y (n_3043));
  NAND3BXL g178543(.AN (n_2601), .B (latched_rd[2]), .C (n_592), .Y
       (n_347));
  NOR3X1 g178544(.A (latched_rd[1]), .B (n_638), .C (n_2598), .Y
       (n_3041));
  OR3X2 g178546(.A (n_580), .B (n_1331), .C (n_2601), .Y (n_3040));
  INVX1 g178547(.A (n_3008), .Y (n_3009));
  INVX1 g178548(.A (n_3005), .Y (n_3006));
  INVX1 g178552(.A (n_2996), .Y (n_2995));
  AOI22X1 g178553(.A0 (\cpuregs[26] [8]), .A1 (n_2493), .B0
       (\cpuregs[28] [8]), .B1 (n_2491), .Y (n_2993));
  AOI22X1 g178554(.A0 (\cpuregs[8] [15]), .A1 (n_2494), .B0
       (\cpuregs[6] [15]), .B1 (n_2530), .Y (n_2992));
  AOI22X1 g178555(.A0 (\cpuregs[9] [15]), .A1 (n_2526), .B0
       (\cpuregs[7] [15]), .B1 (n_12), .Y (n_2991));
  AOI22X1 g178556(.A0 (\cpuregs[10] [15]), .A1 (n_2520), .B0
       (\cpuregs[11] [15]), .B1 (n_2497), .Y (n_2990));
  AOI22X1 g178557(.A0 (\cpuregs[4] [15]), .A1 (n_2529), .B0
       (\cpuregs[5] [15]), .B1 (n_2492), .Y (n_2989));
  AOI22X1 g178558(.A0 (\cpuregs[17] [14]), .A1 (n_2527), .B0
       (\cpuregs[18] [14]), .B1 (n_2519), .Y (n_2988));
  AOI22X1 g178559(.A0 (\cpuregs[20] [14]), .A1 (n_2522), .B0
       (\cpuregs[19] [14]), .B1 (n_2496), .Y (n_2987));
  AOI22X1 g178560(.A0 (\cpuregs[21] [14]), .A1 (n_2495), .B0
       (\cpuregs[22] [14]), .B1 (n_2518), .Y (n_2986));
  AOI22X1 g178561(.A0 (\cpuregs[16] [6]), .A1 (n_2502), .B0
       (\cpuregs[15] [6]), .B1 (n_2504), .Y (n_2985));
  AOI22X1 g178562(.A0 (\cpuregs[26] [14]), .A1 (n_2493), .B0
       (\cpuregs[30] [14]), .B1 (n_2523), .Y (n_2984));
  AOI22X1 g178563(.A0 (\cpuregs[12] [14]), .A1 (n_2521), .B0
       (\cpuregs[13] [14]), .B1 (n_2498), .Y (n_2983));
  AOI22X1 g178564(.A0 (\cpuregs[10] [14]), .A1 (n_2520), .B0
       (\cpuregs[11] [14]), .B1 (n_2497), .Y (n_2982));
  AOI22X1 g178565(.A0 (\cpuregs[2] [14]), .A1 (n_38), .B0
       (\cpuregs[3] [14]), .B1 (n_2503), .Y (n_2981));
  AOI22X1 g178566(.A0 (\cpuregs[4] [14]), .A1 (n_2529), .B0
       (\cpuregs[5] [14]), .B1 (n_2492), .Y (n_2980));
  AOI22X1 g178567(.A0 (\cpuregs[25] [13]), .A1 (n_2528), .B0
       (\cpuregs[26] [13]), .B1 (n_2493), .Y (n_2979));
  AOI22X1 g178568(.A0 (\cpuregs[24] [13]), .A1 (n_2490), .B0
       (\cpuregs[23] [13]), .B1 (n_2500), .Y (n_2978));
  AOI22X1 g178569(.A0 (\cpuregs[29] [13]), .A1 (n_2524), .B0
       (\cpuregs[30] [13]), .B1 (n_2523), .Y (n_2977));
  AOI22X1 g178572(.A0 (\cpuregs[17] [13]), .A1 (n_2527), .B0
       (\cpuregs[20] [13]), .B1 (n_2522), .Y (n_2976));
  AOI22X1 g178573(.A0 (\cpuregs[16] [13]), .A1 (n_2502), .B0
       (\cpuregs[21] [13]), .B1 (n_2495), .Y (n_2975));
  AOI22X1 g178574(.A0 (\cpuregs[19] [13]), .A1 (n_2496), .B0
       (\cpuregs[22] [13]), .B1 (n_2518), .Y (n_2974));
  NOR2X1 g178580(.A (n_544), .B (n_2554), .Y (n_2973));
  NOR2X1 g178581(.A (n_544), .B (n_2566), .Y (n_2972));
  AOI22X1 g178582(.A0 (\cpuregs[8] [13]), .A1 (n_2494), .B0
       (\cpuregs[9] [13]), .B1 (n_2526), .Y (n_2971));
  NOR2X1 g178583(.A (n_544), .B (n_2565), .Y (n_2970));
  NOR2X1 g178584(.A (n_544), .B (n_2553), .Y (n_2969));
  NOR2X1 g178585(.A (n_544), .B (n_2562), .Y (n_2968));
  NOR2X1 g178586(.A (n_2561), .B (n_544), .Y (n_2967));
  NOR2X1 g178587(.A (n_544), .B (n_2552), .Y (n_2966));
  AOI22X1 g178588(.A0 (\cpuregs[6] [13]), .A1 (n_2530), .B0
       (\cpuregs[7] [13]), .B1 (n_12), .Y (n_2965));
  NOR2X1 g178589(.A (n_544), .B (n_2564), .Y (n_2964));
  AOI22X1 g178590(.A0 (\cpuregs[10] [13]), .A1 (n_2520), .B0
       (\cpuregs[11] [13]), .B1 (n_2497), .Y (n_2963));
  AOI22X1 g178591(.A0 (\cpuregs[4] [13]), .A1 (n_2529), .B0
       (\cpuregs[5] [13]), .B1 (n_2492), .Y (n_2962));
  AOI22X1 g178592(.A0 (\cpuregs[17] [12]), .A1 (n_2527), .B0
       (\cpuregs[18] [12]), .B1 (n_2519), .Y (n_2961));
  AOI22X1 g178593(.A0 (\cpuregs[16] [12]), .A1 (n_2502), .B0
       (\cpuregs[15] [12]), .B1 (n_2504), .Y (n_2960));
  AOI22X1 g178594(.A0 (\cpuregs[20] [12]), .A1 (n_2522), .B0
       (\cpuregs[19] [12]), .B1 (n_2496), .Y (n_2959));
  AOI22X1 g178595(.A0 (\cpuregs[24] [7]), .A1 (n_2490), .B0
       (\cpuregs[23] [7]), .B1 (n_2500), .Y (n_2958));
  AOI22X1 g178596(.A0 (\cpuregs[24] [12]), .A1 (n_2490), .B0
       (\cpuregs[23] [12]), .B1 (n_2500), .Y (n_2957));
  AOI22X1 g178597(.A0 (\cpuregs[27] [12]), .A1 (n_2525), .B0
       (\cpuregs[30] [12]), .B1 (n_2523), .Y (n_2956));
  NOR2X1 g178598(.A (n_2434), .B (n_429), .Y (n_2955));
  AOI22X1 g178599(.A0 (\cpuregs[8] [12]), .A1 (n_2494), .B0
       (\cpuregs[6] [12]), .B1 (n_2530), .Y (n_2954));
  AOI22X1 g178600(.A0 (\cpuregs[9] [12]), .A1 (n_2526), .B0
       (\cpuregs[7] [12]), .B1 (n_12), .Y (n_2953));
  AOI22X1 g178601(.A0 (\cpuregs[10] [12]), .A1 (n_2520), .B0
       (\cpuregs[11] [12]), .B1 (n_2497), .Y (n_2952));
  AOI22X1 g178602(.A0 (\cpuregs[12] [12]), .A1 (n_2521), .B0
       (\cpuregs[13] [12]), .B1 (n_2498), .Y (n_2951));
  AOI21X1 g178603(.A0 (n_781), .A1 (n_2483), .B0 (n_544), .Y (n_2950));
  NAND3X1 g178604(.A (n_2045), .B (n_2044), .C (n_2557), .Y (n_2949));
  NAND3X1 g178605(.A (n_2037), .B (n_2036), .C (n_2556), .Y (n_2948));
  NAND4XL g178606(.A (n_542), .B (n_1871), .C (n_2414), .D (n_1632), .Y
       (n_2947));
  AOI22X1 g178607(.A0 (\cpuregs[2] [12]), .A1 (n_38), .B0
       (\cpuregs[3] [12]), .B1 (n_2503), .Y (n_2946));
  AOI22X1 g178608(.A0 (\cpuregs[4] [12]), .A1 (n_2529), .B0
       (\cpuregs[5] [12]), .B1 (n_2492), .Y (n_2945));
  AOI32X1 g178609(.A0 (mem_rdata_q[12]), .A1 (n_538), .A2 (n_2427), .B0
       (instr_sltu), .B1 (n_537), .Y (n_2944));
  NOR4BBX1 g178610(.AN (n_973), .BN (n_2334), .C (n_1638), .D (n_2508),
       .Y (n_2943));
  AOI22X1 g178611(.A0 (\cpuregs[13] [17]), .A1 (n_2498), .B0
       (\cpuregs[7] [17]), .B1 (n_12), .Y (n_2942));
  AOI22X1 g178612(.A0 (\cpuregs[16] [5]), .A1 (n_2502), .B0
       (\cpuregs[15] [5]), .B1 (n_2504), .Y (n_2941));
  AOI22X1 g178613(.A0 (\cpuregs[6] [5]), .A1 (n_2530), .B0
       (\cpuregs[7] [5]), .B1 (n_12), .Y (n_2940));
  AOI22X1 g178614(.A0 (\cpuregs[24] [16]), .A1 (n_2490), .B0
       (\cpuregs[23] [16]), .B1 (n_2500), .Y (n_2939));
  AOI22X1 g178615(.A0 (\cpuregs[28] [16]), .A1 (n_2491), .B0
       (\cpuregs[27] [16]), .B1 (n_2525), .Y (n_2938));
  AOI22X1 g178616(.A0 (\cpuregs[19] [16]), .A1 (n_2496), .B0
       (\cpuregs[22] [16]), .B1 (n_2518), .Y (n_2937));
  AOI22X1 g178617(.A0 (\cpuregs[16] [16]), .A1 (n_2502), .B0
       (\cpuregs[17] [16]), .B1 (n_2527), .Y (n_2936));
  AOI22X1 g178618(.A0 (\cpuregs[29] [5]), .A1 (n_2524), .B0
       (\cpuregs[30] [5]), .B1 (n_2523), .Y (n_2935));
  AOI22X1 g178619(.A0 (\cpuregs[21] [15]), .A1 (n_2495), .B0
       (\cpuregs[22] [15]), .B1 (n_2518), .Y (n_2934));
  AOI22X1 g178620(.A0 (\cpuregs[20] [15]), .A1 (n_2522), .B0
       (\cpuregs[19] [15]), .B1 (n_2496), .Y (n_2933));
  AOI22X1 g178621(.A0 (\cpuregs[17] [28]), .A1 (n_2527), .B0
       (\cpuregs[18] [28]), .B1 (n_2519), .Y (n_2932));
  AOI22X1 g178622(.A0 (\cpuregs[12] [15]), .A1 (n_2521), .B0
       (\cpuregs[13] [15]), .B1 (n_2498), .Y (n_2931));
  AOI22X1 g178623(.A0 (\cpuregs[13] [31]), .A1 (n_2498), .B0
       (\cpuregs[7] [31]), .B1 (n_12), .Y (n_2930));
  AOI22X1 g178624(.A0 (\cpuregs[13] [23]), .A1 (n_2498), .B0
       (\cpuregs[7] [23]), .B1 (n_12), .Y (n_2929));
  AOI22X1 g178625(.A0 (\cpuregs[20] [23]), .A1 (n_2522), .B0
       (\cpuregs[19] [23]), .B1 (n_2496), .Y (n_2928));
  AOI22X1 g178626(.A0 (\cpuregs[17] [10]), .A1 (n_2527), .B0
       (\cpuregs[18] [10]), .B1 (n_2519), .Y (n_2927));
  AOI22X1 g178627(.A0 (\cpuregs[2] [15]), .A1 (n_38), .B0
       (\cpuregs[3] [15]), .B1 (n_2503), .Y (n_2926));
  AOI22X1 g178628(.A0 (\cpuregs[16] [14]), .A1 (n_2502), .B0
       (\cpuregs[15] [14]), .B1 (n_2504), .Y (n_2925));
  AOI22X1 g178629(.A0 (\cpuregs[29] [14]), .A1 (n_2524), .B0
       (\cpuregs[23] [14]), .B1 (n_2500), .Y (n_2924));
  AOI22X1 g178630(.A0 (\cpuregs[25] [14]), .A1 (n_2528), .B0
       (\cpuregs[27] [14]), .B1 (n_2525), .Y (n_2923));
  AOI22X1 g178631(.A0 (\cpuregs[8] [14]), .A1 (n_2494), .B0
       (\cpuregs[9] [14]), .B1 (n_2526), .Y (n_2922));
  AOI22X1 g178632(.A0 (\cpuregs[6] [14]), .A1 (n_2530), .B0
       (\cpuregs[7] [14]), .B1 (n_12), .Y (n_2921));
  AOI22X1 g178633(.A0 (\cpuregs[28] [13]), .A1 (n_2491), .B0
       (\cpuregs[27] [13]), .B1 (n_2525), .Y (n_2920));
  AOI22X1 g178634(.A0 (\cpuregs[4] [5]), .A1 (n_2529), .B0
       (\cpuregs[3] [5]), .B1 (n_2503), .Y (n_2919));
  AOI22X1 g178635(.A0 (\cpuregs[12] [13]), .A1 (n_2521), .B0
       (\cpuregs[13] [13]), .B1 (n_2498), .Y (n_2918));
  AOI22X1 g178636(.A0 (\cpuregs[2] [13]), .A1 (n_38), .B0
       (\cpuregs[3] [13]), .B1 (n_2503), .Y (n_2917));
  AOI22X1 g178637(.A0 (\cpuregs[12] [21]), .A1 (n_2521), .B0
       (\cpuregs[13] [21]), .B1 (n_2498), .Y (n_2916));
  AOI22X1 g178638(.A0 (\cpuregs[21] [12]), .A1 (n_2495), .B0
       (\cpuregs[22] [12]), .B1 (n_2518), .Y (n_2915));
  AOI22X1 g178639(.A0 (\cpuregs[25] [12]), .A1 (n_2528), .B0
       (\cpuregs[29] [12]), .B1 (n_2524), .Y (n_2914));
  AOI22X1 g178640(.A0 (\cpuregs[21] [29]), .A1 (n_2495), .B0
       (\cpuregs[22] [29]), .B1 (n_2518), .Y (n_2913));
  AOI22X1 g178641(.A0 (\cpuregs[5] [10]), .A1 (n_2492), .B0
       (\cpuregs[14] [10]), .B1 (n_2531), .Y (n_2912));
  AOI22X1 g178642(.A0 (\cpuregs[6] [19]), .A1 (n_2530), .B0
       (\cpuregs[7] [19]), .B1 (n_12), .Y (n_2911));
  AOI22X1 g178643(.A0 (\cpuregs[20] [8]), .A1 (n_2522), .B0
       (\cpuregs[19] [8]), .B1 (n_2496), .Y (n_2910));
  AOI22X1 g178644(.A0 (\cpuregs[16] [11]), .A1 (n_2502), .B0
       (\cpuregs[15] [11]), .B1 (n_2504), .Y (n_2909));
  AOI22X1 g178645(.A0 (\cpuregs[21] [11]), .A1 (n_2495), .B0
       (\cpuregs[22] [11]), .B1 (n_2518), .Y (n_2908));
  AOI22X1 g178646(.A0 (\cpuregs[6] [10]), .A1 (n_2530), .B0
       (\cpuregs[7] [10]), .B1 (n_12), .Y (n_2907));
  AOI22X1 g178647(.A0 (\cpuregs[29] [11]), .A1 (n_2524), .B0
       (\cpuregs[23] [11]), .B1 (n_2500), .Y (n_2906));
  AOI22X1 g178648(.A0 (\cpuregs[13] [11]), .A1 (n_2498), .B0
       (\cpuregs[7] [11]), .B1 (n_12), .Y (n_2905));
  AOI22X1 g178649(.A0 (\cpuregs[4] [11]), .A1 (n_2529), .B0
       (\cpuregs[5] [11]), .B1 (n_2492), .Y (n_2904));
  AOI22X1 g178650(.A0 (\cpuregs[2] [11]), .A1 (n_38), .B0
       (\cpuregs[3] [11]), .B1 (n_2503), .Y (n_2903));
  AOI22X1 g178651(.A0 (\cpuregs[16] [10]), .A1 (n_2502), .B0
       (\cpuregs[15] [10]), .B1 (n_2504), .Y (n_2902));
  AOI22X1 g178652(.A0 (\cpuregs[29] [10]), .A1 (n_2524), .B0
       (\cpuregs[30] [10]), .B1 (n_2523), .Y (n_2901));
  AOI22X1 g178653(.A0 (\cpuregs[10] [9]), .A1 (n_2520), .B0
       (\cpuregs[6] [9]), .B1 (n_2530), .Y (n_2900));
  AOI22X1 g178654(.A0 (\cpuregs[6] [27]), .A1 (n_2530), .B0
       (\cpuregs[7] [27]), .B1 (n_12), .Y (n_2899));
  AOI22X1 g178655(.A0 (\cpuregs[8] [10]), .A1 (n_2494), .B0
       (\cpuregs[9] [10]), .B1 (n_2526), .Y (n_2898));
  AOI22X1 g178656(.A0 (\cpuregs[2] [9]), .A1 (n_38), .B0
       (\cpuregs[3] [9]), .B1 (n_2503), .Y (n_2897));
  AOI22X1 g178657(.A0 (\cpuregs[29] [17]), .A1 (n_2524), .B0
       (\cpuregs[30] [17]), .B1 (n_2523), .Y (n_2896));
  AOI22X1 g178658(.A0 (\cpuregs[11] [9]), .A1 (n_2497), .B0
       (\cpuregs[7] [9]), .B1 (n_12), .Y (n_2895));
  AOI22X1 g178659(.A0 (\cpuregs[16] [8]), .A1 (n_2502), .B0
       (\cpuregs[15] [8]), .B1 (n_2504), .Y (n_2894));
  AOI22X1 g178660(.A0 (\cpuregs[17] [11]), .A1 (n_2527), .B0
       (\cpuregs[18] [11]), .B1 (n_2519), .Y (n_2893));
  AOI22X1 g178661(.A0 (\cpuregs[13] [8]), .A1 (n_2498), .B0
       (\cpuregs[7] [8]), .B1 (n_12), .Y (n_2892));
  AOI22X1 g178662(.A0 (\cpuregs[5] [5]), .A1 (n_2492), .B0
       (\cpuregs[14] [5]), .B1 (n_2531), .Y (n_2891));
  AO22X1 g178663(.A0 (\cpuregs[2] [5]), .A1 (n_38), .B0
       (decoded_imm[5]), .B1 (n_421), .Y (n_2890));
  AOI22X1 g178664(.A0 (\cpuregs[12] [5]), .A1 (n_2521), .B0
       (\cpuregs[13] [5]), .B1 (n_2498), .Y (n_2889));
  AOI22X1 g178665(.A0 (\cpuregs[10] [5]), .A1 (n_2520), .B0
       (\cpuregs[11] [5]), .B1 (n_2497), .Y (n_2888));
  AOI22X1 g178666(.A0 (\cpuregs[4] [8]), .A1 (n_2529), .B0
       (\cpuregs[5] [8]), .B1 (n_2492), .Y (n_2887));
  AOI22X1 g178667(.A0 (\cpuregs[8] [5]), .A1 (n_2494), .B0
       (\cpuregs[9] [5]), .B1 (n_2526), .Y (n_2886));
  AOI22X1 g178668(.A0 (\cpuregs[25] [5]), .A1 (n_2528), .B0
       (\cpuregs[26] [5]), .B1 (n_2493), .Y (n_2885));
  AOI22X1 g178669(.A0 (\cpuregs[28] [5]), .A1 (n_2491), .B0
       (\cpuregs[27] [5]), .B1 (n_2525), .Y (n_2884));
  AOI22X1 g178670(.A0 (\cpuregs[24] [5]), .A1 (n_2490), .B0
       (\cpuregs[23] [5]), .B1 (n_2500), .Y (n_2883));
  AOI22X1 g178671(.A0 (\cpuregs[21] [5]), .A1 (n_2495), .B0
       (\cpuregs[22] [5]), .B1 (n_2518), .Y (n_2882));
  AOI22X1 g178672(.A0 (\cpuregs[10] [7]), .A1 (n_2520), .B0
       (\reg_op2[7]_9676 ), .B1 (n_832), .Y (n_2881));
  AOI22X1 g178673(.A0 (\cpuregs[20] [5]), .A1 (n_2522), .B0
       (\cpuregs[19] [5]), .B1 (n_2496), .Y (n_2880));
  AOI22X1 g178674(.A0 (\cpuregs[17] [5]), .A1 (n_2527), .B0
       (\cpuregs[18] [5]), .B1 (n_2519), .Y (n_2879));
  AOI22X1 g178675(.A0 (\cpuregs[5] [6]), .A1 (n_2492), .B0
       (\cpuregs[14] [6]), .B1 (n_2531), .Y (n_2878));
  AOI22X1 g178676(.A0 (\cpuregs[4] [6]), .A1 (n_2529), .B0
       (\cpuregs[3] [6]), .B1 (n_2503), .Y (n_2877));
  AO22X1 g178677(.A0 (\cpuregs[2] [6]), .A1 (n_38), .B0
       (decoded_imm[6]), .B1 (n_421), .Y (n_2876));
  AOI22X1 g178678(.A0 (\cpuregs[10] [6]), .A1 (n_2520), .B0
       (\cpuregs[11] [6]), .B1 (n_2497), .Y (n_2875));
  AOI22X1 g178679(.A0 (\cpuregs[8] [6]), .A1 (n_2494), .B0
       (\cpuregs[9] [6]), .B1 (n_2526), .Y (n_2874));
  AOI22X1 g178680(.A0 (\cpuregs[28] [6]), .A1 (n_2491), .B0
       (\cpuregs[27] [6]), .B1 (n_2525), .Y (n_2873));
  AOI22X1 g178681(.A0 (\cpuregs[25] [6]), .A1 (n_2528), .B0
       (\cpuregs[26] [6]), .B1 (n_2493), .Y (n_2872));
  AOI22X1 g178682(.A0 (\cpuregs[24] [6]), .A1 (n_2490), .B0
       (\cpuregs[23] [6]), .B1 (n_2500), .Y (n_2871));
  AOI22X1 g178683(.A0 (\cpuregs[21] [6]), .A1 (n_2495), .B0
       (\cpuregs[22] [6]), .B1 (n_2518), .Y (n_2870));
  AOI22X1 g178684(.A0 (\cpuregs[20] [6]), .A1 (n_2522), .B0
       (\cpuregs[19] [6]), .B1 (n_2496), .Y (n_2869));
  AOI22X1 g178685(.A0 (\cpuregs[17] [6]), .A1 (n_2527), .B0
       (\cpuregs[18] [6]), .B1 (n_2519), .Y (n_2868));
  AOI22X1 g178686(.A0 (\cpuregs[25] [7]), .A1 (n_2528), .B0
       (\cpuregs[26] [7]), .B1 (n_2493), .Y (n_2867));
  AOI22X1 g178687(.A0 (\cpuregs[28] [7]), .A1 (n_2491), .B0
       (\cpuregs[27] [7]), .B1 (n_2525), .Y (n_2866));
  AOI22X1 g178688(.A0 (\cpuregs[12] [26]), .A1 (n_2521), .B0
       (\cpuregs[13] [26]), .B1 (n_2498), .Y (n_2865));
  AOI22X1 g178689(.A0 (\cpuregs[21] [24]), .A1 (n_2495), .B0
       (\cpuregs[22] [24]), .B1 (n_2518), .Y (n_2864));
  AOI22X1 g178690(.A0 (\cpuregs[2] [7]), .A1 (n_38), .B0
       (\cpuregs[31] [7]), .B1 (n_2499), .Y (n_2863));
  AOI22X1 g178691(.A0 (\cpuregs[4] [7]), .A1 (n_2529), .B0
       (\cpuregs[5] [7]), .B1 (n_2492), .Y (n_2862));
  AOI22X1 g178692(.A0 (\cpuregs[20] [7]), .A1 (n_2522), .B0
       (\cpuregs[19] [7]), .B1 (n_2496), .Y (n_2861));
  AOI22X1 g178693(.A0 (\cpuregs[16] [7]), .A1 (n_2502), .B0
       (\cpuregs[15] [7]), .B1 (n_2504), .Y (n_2860));
  AOI22X1 g178694(.A0 (\cpuregs[21] [7]), .A1 (n_2495), .B0
       (\cpuregs[22] [7]), .B1 (n_2518), .Y (n_2859));
  AOI22X1 g178695(.A0 (\cpuregs[17] [7]), .A1 (n_2527), .B0
       (\cpuregs[18] [7]), .B1 (n_2519), .Y (n_2858));
  AO22X1 g178696(.A0 (\cpuregs[6] [7]), .A1 (n_2530), .B0
       (\cpuregs[13] [7]), .B1 (n_2498), .Y (n_2857));
  AOI22X1 g178697(.A0 (\cpuregs[12] [7]), .A1 (n_2521), .B0
       (\cpuregs[11] [7]), .B1 (n_2497), .Y (n_2856));
  AOI22X1 g178698(.A0 (\cpuregs[2] [8]), .A1 (n_38), .B0
       (\cpuregs[3] [8]), .B1 (n_2503), .Y (n_2855));
  AOI22X1 g178699(.A0 (\cpuregs[12] [8]), .A1 (n_2521), .B0
       (\cpuregs[6] [8]), .B1 (n_2530), .Y (n_2854));
  AOI22X1 g178700(.A0 (\cpuregs[10] [8]), .A1 (n_2520), .B0
       (\cpuregs[11] [8]), .B1 (n_2497), .Y (n_2853));
  AOI22X1 g178701(.A0 (\cpuregs[8] [8]), .A1 (n_2494), .B0
       (\cpuregs[9] [8]), .B1 (n_2526), .Y (n_2852));
  AOI22X1 g178702(.A0 (\cpuregs[29] [8]), .A1 (n_2524), .B0
       (\cpuregs[23] [8]), .B1 (n_2500), .Y (n_2851));
  AOI22X1 g178703(.A0 (\cpuregs[24] [8]), .A1 (n_2490), .B0
       (\cpuregs[25] [8]), .B1 (n_2528), .Y (n_2850));
  AOI22X1 g178704(.A0 (\cpuregs[21] [8]), .A1 (n_2495), .B0
       (\cpuregs[22] [8]), .B1 (n_2518), .Y (n_2849));
  AOI22X1 g178705(.A0 (\cpuregs[17] [8]), .A1 (n_2527), .B0
       (\cpuregs[18] [8]), .B1 (n_2519), .Y (n_2848));
  AOI22X1 g178706(.A0 (\cpuregs[4] [9]), .A1 (n_2529), .B0
       (\cpuregs[5] [9]), .B1 (n_2492), .Y (n_2847));
  AOI22X1 g178707(.A0 (\cpuregs[12] [9]), .A1 (n_2521), .B0
       (\cpuregs[13] [9]), .B1 (n_2498), .Y (n_2846));
  AOI22X1 g178708(.A0 (\cpuregs[8] [9]), .A1 (n_2494), .B0
       (\cpuregs[9] [9]), .B1 (n_2526), .Y (n_2845));
  AOI22X1 g178709(.A0 (\cpuregs[26] [9]), .A1 (n_2493), .B0
       (\cpuregs[23] [9]), .B1 (n_2500), .Y (n_2844));
  AOI22X1 g178710(.A0 (\cpuregs[25] [9]), .A1 (n_2528), .B0
       (\cpuregs[27] [9]), .B1 (n_2525), .Y (n_2843));
  AOI22X1 g178711(.A0 (\cpuregs[24] [9]), .A1 (n_2490), .B0
       (\cpuregs[30] [9]), .B1 (n_2523), .Y (n_2842));
  AOI22X1 g178712(.A0 (\cpuregs[21] [9]), .A1 (n_2495), .B0
       (\cpuregs[22] [9]), .B1 (n_2518), .Y (n_2841));
  AOI22X1 g178713(.A0 (\cpuregs[16] [9]), .A1 (n_2502), .B0
       (\cpuregs[15] [9]), .B1 (n_2504), .Y (n_2840));
  AOI22X1 g178714(.A0 (\cpuregs[20] [9]), .A1 (n_2522), .B0
       (\cpuregs[19] [9]), .B1 (n_2496), .Y (n_2839));
  AOI22X1 g178715(.A0 (\cpuregs[17] [9]), .A1 (n_2527), .B0
       (\cpuregs[18] [9]), .B1 (n_2519), .Y (n_2838));
  AOI22X1 g178716(.A0 (\cpuregs[4] [10]), .A1 (n_2529), .B0
       (\cpuregs[3] [10]), .B1 (n_2503), .Y (n_2837));
  AO22X1 g178717(.A0 (\cpuregs[2] [10]), .A1 (n_38), .B0
       (decoded_imm[10]), .B1 (n_421), .Y (n_2836));
  AOI22X1 g178718(.A0 (\cpuregs[12] [10]), .A1 (n_2521), .B0
       (\cpuregs[13] [10]), .B1 (n_2498), .Y (n_2835));
  AOI22X1 g178719(.A0 (\cpuregs[10] [10]), .A1 (n_2520), .B0
       (\cpuregs[11] [10]), .B1 (n_2497), .Y (n_2834));
  AOI22X1 g178720(.A0 (\cpuregs[25] [10]), .A1 (n_2528), .B0
       (\cpuregs[26] [10]), .B1 (n_2493), .Y (n_2833));
  AOI22X1 g178721(.A0 (\cpuregs[28] [10]), .A1 (n_2491), .B0
       (\cpuregs[23] [10]), .B1 (n_2500), .Y (n_2832));
  AOI22X1 g178722(.A0 (\cpuregs[24] [10]), .A1 (n_2490), .B0
       (\cpuregs[27] [10]), .B1 (n_2525), .Y (n_2831));
  AOI22X1 g178723(.A0 (\cpuregs[21] [10]), .A1 (n_2495), .B0
       (\cpuregs[22] [10]), .B1 (n_2518), .Y (n_2830));
  AOI22X1 g178724(.A0 (\cpuregs[20] [10]), .A1 (n_2522), .B0
       (\cpuregs[19] [10]), .B1 (n_2496), .Y (n_2829));
  AOI22X1 g178725(.A0 (\cpuregs[12] [11]), .A1 (n_2521), .B0
       (\cpuregs[6] [11]), .B1 (n_2530), .Y (n_2828));
  AOI22X1 g178726(.A0 (\cpuregs[10] [11]), .A1 (n_2520), .B0
       (\cpuregs[11] [11]), .B1 (n_2497), .Y (n_2827));
  AOI22X1 g178727(.A0 (\cpuregs[8] [11]), .A1 (n_2494), .B0
       (\cpuregs[9] [11]), .B1 (n_2526), .Y (n_2826));
  AOI22X1 g178728(.A0 (\cpuregs[24] [11]), .A1 (n_2490), .B0
       (\cpuregs[28] [11]), .B1 (n_2491), .Y (n_2825));
  AOI22X1 g178729(.A0 (\cpuregs[25] [11]), .A1 (n_2528), .B0
       (\cpuregs[27] [11]), .B1 (n_2525), .Y (n_2824));
  AOI22X1 g178730(.A0 (\cpuregs[20] [11]), .A1 (n_2522), .B0
       (\cpuregs[19] [11]), .B1 (n_2496), .Y (n_2823));
  NAND2BX1 g178735(.AN (n_429), .B (n_13), .Y (n_3008));
  AOI21X1 g178736(.A0 (n_2515), .A1 (n_1589), .B0 (n_2421), .Y
       (n_3007));
  AOI21X1 g178737(.A0 (n_2514), .A1 (n_2433), .B0 (n_2506), .Y
       (n_3005));
  NOR2X1 g178739(.A (n_592), .B (n_2598), .Y (n_3004));
  NOR2X1 g178741(.A (decoded_rs1[3]), .B (n_2586), .Y (n_3003));
  NAND2BX1 g178742(.AN (n_2586), .B (decoded_rs1[3]), .Y (n_3002));
  NOR2X1 g178743(.A (n_592), .B (n_2601), .Y (n_3001));
  NOR2BX1 g178744(.AN (n_979), .B (n_2601), .Y (n_3000));
  NOR2BX1 g178745(.AN (n_979), .B (n_2598), .Y (n_2999));
  AND2X1 g178762(.A (n_1589), .B (n_2599), .Y (n_2998));
  NOR2X1 g178763(.A (n_2423), .B (n_2607), .Y (n_2997));
  NAND2X1 g178764(.A (n_2131), .B (n_429), .Y (n_2996));
  AND2X2 g178765(.A (n_580), .B (n_11747), .Y (n_508));
  AOI22X1 g178767(.A0 (\cpuregs[20] [24]), .A1 (n_2522), .B0
       (\cpuregs[19] [24]), .B1 (n_2496), .Y (n_2821));
  AOI22X1 g178768(.A0 (\cpuregs[24] [15]), .A1 (n_2490), .B0
       (\cpuregs[23] [15]), .B1 (n_2500), .Y (n_2820));
  AOI22X1 g178769(.A0 (\cpuregs[26] [15]), .A1 (n_2493), .B0
       (\cpuregs[30] [15]), .B1 (n_2523), .Y (n_2819));
  AOI22X1 g178770(.A0 (\cpuregs[16] [15]), .A1 (n_2502), .B0
       (\cpuregs[15] [15]), .B1 (n_2504), .Y (n_2818));
  AOI22X1 g178771(.A0 (\cpuregs[17] [15]), .A1 (n_2527), .B0
       (\cpuregs[18] [15]), .B1 (n_2519), .Y (n_2817));
  AOI22X1 g178772(.A0 (\cpuregs[4] [16]), .A1 (n_2529), .B0
       (\cpuregs[5] [16]), .B1 (n_2492), .Y (n_2816));
  AOI22X1 g178773(.A0 (\cpuregs[2] [16]), .A1 (n_38), .B0
       (\cpuregs[3] [16]), .B1 (n_2503), .Y (n_2815));
  AOI22X1 g178774(.A0 (\cpuregs[11] [16]), .A1 (n_2497), .B0
       (\cpuregs[7] [16]), .B1 (n_12), .Y (n_2814));
  AOI22X1 g178775(.A0 (\cpuregs[10] [16]), .A1 (n_2520), .B0
       (\cpuregs[6] [16]), .B1 (n_2530), .Y (n_2813));
  AOI22X1 g178776(.A0 (\cpuregs[12] [16]), .A1 (n_2521), .B0
       (\cpuregs[13] [16]), .B1 (n_2498), .Y (n_2812));
  AOI22X1 g178777(.A0 (\cpuregs[8] [16]), .A1 (n_2494), .B0
       (\cpuregs[9] [16]), .B1 (n_2526), .Y (n_2811));
  AOI22X1 g178778(.A0 (\cpuregs[18] [16]), .A1 (n_2519), .B0
       (\cpuregs[21] [16]), .B1 (n_2495), .Y (n_2810));
  AOI22X1 g178779(.A0 (\cpuregs[29] [16]), .A1 (n_2524), .B0
       (\cpuregs[30] [16]), .B1 (n_2523), .Y (n_2809));
  AOI22X1 g178780(.A0 (\cpuregs[25] [16]), .A1 (n_2528), .B0
       (\cpuregs[26] [16]), .B1 (n_2493), .Y (n_2808));
  AOI22X1 g178781(.A0 (\cpuregs[5] [17]), .A1 (n_2492), .B0
       (\cpuregs[14] [17]), .B1 (n_2531), .Y (n_2807));
  AOI22X1 g178782(.A0 (\cpuregs[4] [17]), .A1 (n_2529), .B0
       (\cpuregs[3] [17]), .B1 (n_2503), .Y (n_2806));
  AO22X1 g178783(.A0 (\cpuregs[2] [17]), .A1 (n_38), .B0
       (decoded_imm[17]), .B1 (n_421), .Y (n_2805));
  AOI22X1 g178784(.A0 (\cpuregs[12] [17]), .A1 (n_2521), .B0
       (\cpuregs[6] [17]), .B1 (n_2530), .Y (n_2804));
  AOI22X1 g178785(.A0 (\cpuregs[10] [17]), .A1 (n_2520), .B0
       (\cpuregs[11] [17]), .B1 (n_2497), .Y (n_2803));
  AOI22X1 g178786(.A0 (\cpuregs[8] [17]), .A1 (n_2494), .B0
       (\cpuregs[9] [17]), .B1 (n_2526), .Y (n_2802));
  AOI22X1 g178787(.A0 (\cpuregs[25] [17]), .A1 (n_2528), .B0
       (\cpuregs[26] [17]), .B1 (n_2493), .Y (n_2801));
  AOI22X1 g178788(.A0 (\cpuregs[24] [17]), .A1 (n_2490), .B0
       (\cpuregs[23] [17]), .B1 (n_2500), .Y (n_2800));
  AOI22X1 g178789(.A0 (\cpuregs[21] [17]), .A1 (n_2495), .B0
       (\cpuregs[22] [17]), .B1 (n_2518), .Y (n_2799));
  AOI22X1 g178790(.A0 (\cpuregs[16] [17]), .A1 (n_2502), .B0
       (\cpuregs[15] [17]), .B1 (n_2504), .Y (n_2798));
  AOI22X1 g178791(.A0 (\cpuregs[20] [17]), .A1 (n_2522), .B0
       (\cpuregs[19] [17]), .B1 (n_2496), .Y (n_2797));
  AOI22X1 g178792(.A0 (\cpuregs[17] [17]), .A1 (n_2527), .B0
       (\cpuregs[18] [17]), .B1 (n_2519), .Y (n_2796));
  AOI22X1 g178793(.A0 (\cpuregs[4] [18]), .A1 (n_2529), .B0
       (\cpuregs[5] [18]), .B1 (n_2492), .Y (n_2795));
  AOI22X1 g178794(.A0 (\cpuregs[2] [18]), .A1 (n_38), .B0
       (\cpuregs[3] [18]), .B1 (n_2503), .Y (n_2794));
  AOI22X1 g178795(.A0 (\cpuregs[6] [18]), .A1 (n_2530), .B0
       (\cpuregs[7] [18]), .B1 (n_12), .Y (n_2793));
  AOI22X1 g178796(.A0 (\cpuregs[10] [18]), .A1 (n_2520), .B0
       (\cpuregs[11] [18]), .B1 (n_2497), .Y (n_2792));
  AOI22X1 g178797(.A0 (\cpuregs[12] [18]), .A1 (n_2521), .B0
       (\cpuregs[13] [18]), .B1 (n_2498), .Y (n_2791));
  AOI22X1 g178798(.A0 (\cpuregs[8] [18]), .A1 (n_2494), .B0
       (\cpuregs[9] [18]), .B1 (n_2526), .Y (n_2790));
  AOI22X1 g178799(.A0 (\cpuregs[27] [18]), .A1 (n_2525), .B0
       (\cpuregs[30] [18]), .B1 (n_2523), .Y (n_2789));
  AOI22X1 g178800(.A0 (\cpuregs[24] [18]), .A1 (n_2490), .B0
       (\cpuregs[23] [18]), .B1 (n_2500), .Y (n_2788));
  AOI22X1 g178801(.A0 (\cpuregs[25] [18]), .A1 (n_2528), .B0
       (\cpuregs[29] [18]), .B1 (n_2524), .Y (n_2787));
  AOI22X1 g178802(.A0 (\cpuregs[29] [6]), .A1 (n_2524), .B0
       (\cpuregs[30] [6]), .B1 (n_2523), .Y (n_2786));
  AOI22X1 g178803(.A0 (\cpuregs[21] [18]), .A1 (n_2495), .B0
       (\cpuregs[22] [18]), .B1 (n_2518), .Y (n_2785));
  AOI22X1 g178804(.A0 (\cpuregs[20] [18]), .A1 (n_2522), .B0
       (\cpuregs[19] [18]), .B1 (n_2496), .Y (n_2784));
  AOI22X1 g178805(.A0 (\cpuregs[16] [18]), .A1 (n_2502), .B0
       (\cpuregs[15] [18]), .B1 (n_2504), .Y (n_2783));
  AOI22X1 g178806(.A0 (\cpuregs[17] [18]), .A1 (n_2527), .B0
       (\cpuregs[18] [18]), .B1 (n_2519), .Y (n_2782));
  AOI22X1 g178807(.A0 (\cpuregs[4] [19]), .A1 (n_2529), .B0
       (\cpuregs[5] [19]), .B1 (n_2492), .Y (n_2781));
  AOI22X1 g178808(.A0 (\cpuregs[2] [19]), .A1 (n_38), .B0
       (\cpuregs[3] [19]), .B1 (n_2503), .Y (n_2780));
  AOI22X1 g178809(.A0 (\cpuregs[12] [19]), .A1 (n_2521), .B0
       (\cpuregs[13] [19]), .B1 (n_2498), .Y (n_2779));
  AOI22X1 g178810(.A0 (\cpuregs[10] [19]), .A1 (n_2520), .B0
       (\cpuregs[11] [19]), .B1 (n_2497), .Y (n_2778));
  AOI22X1 g178811(.A0 (\cpuregs[8] [19]), .A1 (n_2494), .B0
       (\cpuregs[9] [19]), .B1 (n_2526), .Y (n_2777));
  AOI22X1 g178812(.A0 (\cpuregs[27] [19]), .A1 (n_2525), .B0
       (\cpuregs[23] [19]), .B1 (n_2500), .Y (n_2776));
  AOI22X1 g178813(.A0 (\cpuregs[28] [19]), .A1 (n_2491), .B0
       (\cpuregs[29] [19]), .B1 (n_2524), .Y (n_2775));
  AOI22X1 g178814(.A0 (\cpuregs[24] [19]), .A1 (n_2490), .B0
       (\cpuregs[25] [19]), .B1 (n_2528), .Y (n_2774));
  AOI22X1 g178815(.A0 (\cpuregs[20] [19]), .A1 (n_2522), .B0
       (\cpuregs[19] [19]), .B1 (n_2496), .Y (n_2773));
  AOI22X1 g178816(.A0 (\cpuregs[16] [19]), .A1 (n_2502), .B0
       (\cpuregs[15] [19]), .B1 (n_2504), .Y (n_2772));
  AOI22X1 g178817(.A0 (\cpuregs[21] [19]), .A1 (n_2495), .B0
       (\cpuregs[22] [19]), .B1 (n_2518), .Y (n_2771));
  AOI22X1 g178818(.A0 (\cpuregs[17] [19]), .A1 (n_2527), .B0
       (\cpuregs[18] [19]), .B1 (n_2519), .Y (n_2770));
  AOI22X1 g178819(.A0 (\cpuregs[4] [20]), .A1 (n_2529), .B0
       (\cpuregs[5] [20]), .B1 (n_2492), .Y (n_2769));
  AOI22X1 g178820(.A0 (\cpuregs[2] [20]), .A1 (n_38), .B0
       (\cpuregs[3] [20]), .B1 (n_2503), .Y (n_2768));
  AOI22X1 g178821(.A0 (\cpuregs[12] [20]), .A1 (n_2521), .B0
       (\cpuregs[13] [20]), .B1 (n_2498), .Y (n_2767));
  AOI22X1 g178822(.A0 (\cpuregs[10] [20]), .A1 (n_2520), .B0
       (\cpuregs[11] [20]), .B1 (n_2497), .Y (n_2766));
  AOI22X1 g178823(.A0 (\cpuregs[6] [20]), .A1 (n_2530), .B0
       (\cpuregs[7] [20]), .B1 (n_12), .Y (n_2765));
  AOI22X1 g178824(.A0 (\cpuregs[8] [20]), .A1 (n_2494), .B0
       (\cpuregs[9] [20]), .B1 (n_2526), .Y (n_2764));
  AOI22X1 g178825(.A0 (\cpuregs[16] [20]), .A1 (n_2502), .B0
       (\cpuregs[19] [20]), .B1 (n_2496), .Y (n_2763));
  AOI22X1 g178826(.A0 (\cpuregs[17] [20]), .A1 (n_2527), .B0
       (\cpuregs[20] [20]), .B1 (n_2522), .Y (n_2762));
  AOI22X1 g178827(.A0 (\cpuregs[18] [20]), .A1 (n_2519), .B0
       (\cpuregs[21] [20]), .B1 (n_2495), .Y (n_2761));
  AOI22X1 g178828(.A0 (\cpuregs[29] [20]), .A1 (n_2524), .B0
       (\cpuregs[30] [20]), .B1 (n_2523), .Y (n_2760));
  AOI22X1 g178829(.A0 (\cpuregs[28] [20]), .A1 (n_2491), .B0
       (\cpuregs[27] [20]), .B1 (n_2525), .Y (n_2759));
  AOI22X1 g178830(.A0 (\cpuregs[25] [20]), .A1 (n_2528), .B0
       (\cpuregs[26] [20]), .B1 (n_2493), .Y (n_2758));
  AOI22X1 g178831(.A0 (\cpuregs[24] [20]), .A1 (n_2490), .B0
       (\cpuregs[23] [20]), .B1 (n_2500), .Y (n_2757));
  AOI22X1 g178832(.A0 (\cpuregs[4] [21]), .A1 (n_2529), .B0
       (\cpuregs[5] [21]), .B1 (n_2492), .Y (n_2756));
  AOI22X1 g178833(.A0 (\cpuregs[2] [21]), .A1 (n_38), .B0
       (\cpuregs[3] [21]), .B1 (n_2503), .Y (n_2755));
  AOI22X1 g178834(.A0 (\cpuregs[10] [21]), .A1 (n_2520), .B0
       (\cpuregs[11] [21]), .B1 (n_2497), .Y (n_2754));
  AOI22X1 g178835(.A0 (\cpuregs[9] [21]), .A1 (n_2526), .B0
       (\cpuregs[7] [21]), .B1 (n_12), .Y (n_2753));
  AOI22X1 g178836(.A0 (\cpuregs[8] [21]), .A1 (n_2494), .B0
       (\cpuregs[6] [21]), .B1 (n_2530), .Y (n_2752));
  AOI22X1 g178837(.A0 (\cpuregs[27] [21]), .A1 (n_2525), .B0
       (\cpuregs[23] [21]), .B1 (n_2500), .Y (n_2751));
  AOI22X1 g178838(.A0 (\cpuregs[28] [21]), .A1 (n_2491), .B0
       (\cpuregs[29] [21]), .B1 (n_2524), .Y (n_2750));
  AOI22X1 g178839(.A0 (\cpuregs[24] [21]), .A1 (n_2490), .B0
       (\cpuregs[25] [21]), .B1 (n_2528), .Y (n_2749));
  AOI22X1 g178840(.A0 (\cpuregs[20] [21]), .A1 (n_2522), .B0
       (\cpuregs[19] [21]), .B1 (n_2496), .Y (n_2748));
  AOI22X1 g178841(.A0 (\cpuregs[16] [21]), .A1 (n_2502), .B0
       (\cpuregs[15] [21]), .B1 (n_2504), .Y (n_2747));
  AOI22X1 g178842(.A0 (\cpuregs[21] [21]), .A1 (n_2495), .B0
       (\cpuregs[22] [21]), .B1 (n_2518), .Y (n_2746));
  AOI22X1 g178843(.A0 (\cpuregs[17] [21]), .A1 (n_2527), .B0
       (\cpuregs[18] [21]), .B1 (n_2519), .Y (n_2745));
  AOI22X1 g178844(.A0 (\cpuregs[4] [22]), .A1 (n_2529), .B0
       (\cpuregs[5] [22]), .B1 (n_2492), .Y (n_2744));
  AOI22X1 g178845(.A0 (\cpuregs[2] [22]), .A1 (n_38), .B0
       (\cpuregs[3] [22]), .B1 (n_2503), .Y (n_2743));
  AOI22X1 g178846(.A0 (\cpuregs[11] [22]), .A1 (n_2497), .B0
       (\cpuregs[7] [22]), .B1 (n_12), .Y (n_2742));
  AOI22X1 g178847(.A0 (\cpuregs[10] [22]), .A1 (n_2520), .B0
       (\cpuregs[6] [22]), .B1 (n_2530), .Y (n_2741));
  AOI22X1 g178848(.A0 (\cpuregs[12] [22]), .A1 (n_2521), .B0
       (\cpuregs[13] [22]), .B1 (n_2498), .Y (n_2740));
  AOI22X1 g178849(.A0 (\cpuregs[8] [22]), .A1 (n_2494), .B0
       (\cpuregs[9] [22]), .B1 (n_2526), .Y (n_2739));
  AOI22X1 g178850(.A0 (\cpuregs[27] [22]), .A1 (n_2525), .B0
       (\cpuregs[30] [22]), .B1 (n_2523), .Y (n_2738));
  AOI22X1 g178851(.A0 (\cpuregs[24] [22]), .A1 (n_2490), .B0
       (\cpuregs[23] [22]), .B1 (n_2500), .Y (n_2737));
  AOI22X1 g178852(.A0 (\cpuregs[25] [22]), .A1 (n_2528), .B0
       (\cpuregs[29] [22]), .B1 (n_2524), .Y (n_2736));
  AOI22X1 g178853(.A0 (\cpuregs[20] [22]), .A1 (n_2522), .B0
       (\cpuregs[19] [22]), .B1 (n_2496), .Y (n_2735));
  AOI22X1 g178854(.A0 (\cpuregs[16] [22]), .A1 (n_2502), .B0
       (\cpuregs[15] [22]), .B1 (n_2504), .Y (n_2734));
  AOI22X1 g178855(.A0 (\cpuregs[21] [22]), .A1 (n_2495), .B0
       (\cpuregs[22] [22]), .B1 (n_2518), .Y (n_2733));
  AOI22X1 g178856(.A0 (\cpuregs[17] [22]), .A1 (n_2527), .B0
       (\cpuregs[18] [22]), .B1 (n_2519), .Y (n_2732));
  AOI22X1 g178857(.A0 (\cpuregs[5] [23]), .A1 (n_2492), .B0
       (\cpuregs[14] [23]), .B1 (n_2531), .Y (n_2731));
  AOI22X1 g178858(.A0 (\cpuregs[4] [23]), .A1 (n_2529), .B0
       (\cpuregs[3] [23]), .B1 (n_2503), .Y (n_2730));
  AO22X1 g178859(.A0 (\cpuregs[2] [23]), .A1 (n_38), .B0
       (decoded_imm[23]), .B1 (n_421), .Y (n_2729));
  AOI22X1 g178860(.A0 (\cpuregs[12] [23]), .A1 (n_2521), .B0
       (\cpuregs[6] [23]), .B1 (n_2530), .Y (n_2728));
  AOI22X1 g178861(.A0 (\cpuregs[10] [23]), .A1 (n_2520), .B0
       (\cpuregs[11] [23]), .B1 (n_2497), .Y (n_2727));
  AOI22X1 g178862(.A0 (\cpuregs[8] [23]), .A1 (n_2494), .B0
       (\cpuregs[9] [23]), .B1 (n_2526), .Y (n_2726));
  AOI22X1 g178863(.A0 (\cpuregs[28] [23]), .A1 (n_2491), .B0
       (\cpuregs[27] [23]), .B1 (n_2525), .Y (n_2725));
  AOI22X1 g178864(.A0 (\cpuregs[25] [23]), .A1 (n_2528), .B0
       (\cpuregs[26] [23]), .B1 (n_2493), .Y (n_2724));
  AOI22X1 g178865(.A0 (\cpuregs[24] [23]), .A1 (n_2490), .B0
       (\cpuregs[23] [23]), .B1 (n_2500), .Y (n_2723));
  AOI22X1 g178866(.A0 (\cpuregs[21] [23]), .A1 (n_2495), .B0
       (\cpuregs[22] [23]), .B1 (n_2518), .Y (n_2722));
  AOI22X1 g178867(.A0 (\cpuregs[16] [23]), .A1 (n_2502), .B0
       (\cpuregs[15] [23]), .B1 (n_2504), .Y (n_2721));
  AOI22X1 g178868(.A0 (\cpuregs[17] [23]), .A1 (n_2527), .B0
       (\cpuregs[18] [23]), .B1 (n_2519), .Y (n_2720));
  AOI22X1 g178869(.A0 (\cpuregs[28] [24]), .A1 (n_2491), .B0
       (\cpuregs[27] [24]), .B1 (n_2525), .Y (n_2719));
  AOI22X1 g178870(.A0 (\cpuregs[25] [24]), .A1 (n_2528), .B0
       (\cpuregs[26] [24]), .B1 (n_2493), .Y (n_2718));
  AOI22X1 g178871(.A0 (\cpuregs[29] [24]), .A1 (n_2524), .B0
       (\cpuregs[30] [24]), .B1 (n_2523), .Y (n_2717));
  AOI22X1 g178872(.A0 (\cpuregs[4] [24]), .A1 (n_2529), .B0
       (\cpuregs[31] [24]), .B1 (n_2499), .Y (n_2716));
  AOI22X1 g178873(.A0 (\cpuregs[2] [24]), .A1 (n_38), .B0
       (\cpuregs[3] [24]), .B1 (n_2503), .Y (n_2715));
  AOI22X1 g178874(.A0 (\cpuregs[25] [15]), .A1 (n_2528), .B0
       (\cpuregs[27] [15]), .B1 (n_2525), .Y (n_2714));
  AOI22X1 g178875(.A0 (\cpuregs[16] [24]), .A1 (n_2502), .B0
       (\cpuregs[15] [24]), .B1 (n_2504), .Y (n_2713));
  AOI22X1 g178876(.A0 (\cpuregs[17] [24]), .A1 (n_2527), .B0
       (\cpuregs[18] [24]), .B1 (n_2519), .Y (n_2712));
  AO22X1 g178877(.A0 (\cpuregs[6] [24]), .A1 (n_2530), .B0
       (\cpuregs[11] [24]), .B1 (n_2497), .Y (n_2711));
  AOI22X1 g178878(.A0 (\cpuregs[8] [24]), .A1 (n_2494), .B0
       (\reg_op2[24]_9693 ), .B1 (n_832), .Y (n_2710));
  AOI22X1 g178879(.A0 (\cpuregs[9] [24]), .A1 (n_2526), .B0
       (\cpuregs[12] [24]), .B1 (n_2521), .Y (n_2709));
  AOI22X1 g178880(.A0 (\cpuregs[2] [25]), .A1 (n_38), .B0
       (\cpuregs[3] [25]), .B1 (n_2503), .Y (n_2708));
  AOI22X1 g178881(.A0 (\cpuregs[4] [25]), .A1 (n_2529), .B0
       (\cpuregs[5] [25]), .B1 (n_2492), .Y (n_2707));
  AOI22X1 g178882(.A0 (\cpuregs[11] [25]), .A1 (n_2497), .B0
       (\cpuregs[7] [25]), .B1 (n_12), .Y (n_2706));
  AOI22X1 g178883(.A0 (\cpuregs[10] [25]), .A1 (n_2520), .B0
       (\cpuregs[6] [25]), .B1 (n_2530), .Y (n_2705));
  AOI22X1 g178884(.A0 (\cpuregs[12] [25]), .A1 (n_2521), .B0
       (\cpuregs[13] [25]), .B1 (n_2498), .Y (n_2704));
  AOI22X1 g178885(.A0 (\cpuregs[8] [25]), .A1 (n_2494), .B0
       (\cpuregs[9] [25]), .B1 (n_2526), .Y (n_2703));
  AOI22X1 g178886(.A0 (\cpuregs[29] [25]), .A1 (n_2524), .B0
       (\cpuregs[23] [25]), .B1 (n_2500), .Y (n_2702));
  AOI22X1 g178887(.A0 (\cpuregs[24] [25]), .A1 (n_2490), .B0
       (\cpuregs[25] [25]), .B1 (n_2528), .Y (n_2701));
  AOI22X1 g178888(.A0 (\cpuregs[26] [25]), .A1 (n_2493), .B0
       (\cpuregs[28] [25]), .B1 (n_2491), .Y (n_2700));
  AOI22X1 g178889(.A0 (\cpuregs[21] [25]), .A1 (n_2495), .B0
       (\cpuregs[22] [25]), .B1 (n_2518), .Y (n_2699));
  AOI22X1 g178890(.A0 (\cpuregs[16] [25]), .A1 (n_2502), .B0
       (\cpuregs[15] [25]), .B1 (n_2504), .Y (n_2698));
  AOI22X1 g178891(.A0 (\cpuregs[20] [25]), .A1 (n_2522), .B0
       (\cpuregs[19] [25]), .B1 (n_2496), .Y (n_2697));
  AOI22X1 g178892(.A0 (\cpuregs[17] [25]), .A1 (n_2527), .B0
       (\cpuregs[18] [25]), .B1 (n_2519), .Y (n_2696));
  AOI22X1 g178893(.A0 (\cpuregs[5] [26]), .A1 (n_2492), .B0
       (\cpuregs[14] [26]), .B1 (n_2531), .Y (n_2695));
  AOI22X1 g178894(.A0 (\cpuregs[4] [26]), .A1 (n_2529), .B0
       (\cpuregs[3] [26]), .B1 (n_2503), .Y (n_2694));
  AO22X1 g178895(.A0 (\cpuregs[2] [26]), .A1 (n_38), .B0
       (decoded_imm[26]), .B1 (n_421), .Y (n_2693));
  AOI22X1 g178896(.A0 (\cpuregs[10] [26]), .A1 (n_2520), .B0
       (\cpuregs[11] [26]), .B1 (n_2497), .Y (n_2692));
  AOI22X1 g178897(.A0 (\cpuregs[6] [26]), .A1 (n_2530), .B0
       (\cpuregs[7] [26]), .B1 (n_12), .Y (n_2691));
  AOI22X1 g178898(.A0 (\cpuregs[8] [26]), .A1 (n_2494), .B0
       (\cpuregs[9] [26]), .B1 (n_2526), .Y (n_2690));
  AOI22X1 g178899(.A0 (\cpuregs[29] [26]), .A1 (n_2524), .B0
       (\cpuregs[30] [26]), .B1 (n_2523), .Y (n_2689));
  AOI22X1 g178900(.A0 (\cpuregs[24] [26]), .A1 (n_2490), .B0
       (\cpuregs[23] [26]), .B1 (n_2500), .Y (n_2688));
  AOI22X1 g178901(.A0 (\cpuregs[28] [26]), .A1 (n_2491), .B0
       (\cpuregs[27] [26]), .B1 (n_2525), .Y (n_2687));
  AOI22X1 g178902(.A0 (\cpuregs[25] [26]), .A1 (n_2528), .B0
       (\cpuregs[26] [26]), .B1 (n_2493), .Y (n_2686));
  AOI22X1 g178903(.A0 (\cpuregs[21] [26]), .A1 (n_2495), .B0
       (\cpuregs[22] [26]), .B1 (n_2518), .Y (n_2685));
  AOI22X1 g178904(.A0 (\cpuregs[20] [26]), .A1 (n_2522), .B0
       (\cpuregs[19] [26]), .B1 (n_2496), .Y (n_2684));
  AOI22X1 g178905(.A0 (\cpuregs[16] [26]), .A1 (n_2502), .B0
       (\cpuregs[15] [26]), .B1 (n_2504), .Y (n_2683));
  AOI22X1 g178906(.A0 (\cpuregs[17] [26]), .A1 (n_2527), .B0
       (\cpuregs[18] [26]), .B1 (n_2519), .Y (n_2682));
  AOI22X1 g178907(.A0 (\cpuregs[4] [27]), .A1 (n_2529), .B0
       (\cpuregs[5] [27]), .B1 (n_2492), .Y (n_2681));
  AOI22X1 g178908(.A0 (\cpuregs[2] [27]), .A1 (n_38), .B0
       (\cpuregs[3] [27]), .B1 (n_2503), .Y (n_2680));
  AOI22X1 g178909(.A0 (\cpuregs[12] [27]), .A1 (n_2521), .B0
       (\cpuregs[13] [27]), .B1 (n_2498), .Y (n_2679));
  AOI22X1 g178910(.A0 (\cpuregs[10] [27]), .A1 (n_2520), .B0
       (\cpuregs[11] [27]), .B1 (n_2497), .Y (n_2678));
  AOI22X1 g178911(.A0 (\cpuregs[8] [27]), .A1 (n_2494), .B0
       (\cpuregs[9] [27]), .B1 (n_2526), .Y (n_2677));
  AOI22X1 g178912(.A0 (\cpuregs[29] [27]), .A1 (n_2524), .B0
       (\cpuregs[23] [27]), .B1 (n_2500), .Y (n_2676));
  AOI22X1 g178913(.A0 (\cpuregs[24] [27]), .A1 (n_2490), .B0
       (\cpuregs[25] [27]), .B1 (n_2528), .Y (n_2675));
  AOI22X1 g178914(.A0 (\cpuregs[26] [27]), .A1 (n_2493), .B0
       (\cpuregs[28] [27]), .B1 (n_2491), .Y (n_2674));
  AOI22X1 g178915(.A0 (\cpuregs[21] [27]), .A1 (n_2495), .B0
       (\cpuregs[22] [27]), .B1 (n_2518), .Y (n_2673));
  AOI22X1 g178916(.A0 (\cpuregs[16] [27]), .A1 (n_2502), .B0
       (\cpuregs[15] [27]), .B1 (n_2504), .Y (n_2672));
  AOI22X1 g178917(.A0 (\cpuregs[20] [27]), .A1 (n_2522), .B0
       (\cpuregs[19] [27]), .B1 (n_2496), .Y (n_2671));
  AOI22X1 g178918(.A0 (\cpuregs[17] [27]), .A1 (n_2527), .B0
       (\cpuregs[18] [27]), .B1 (n_2519), .Y (n_2670));
  AOI22X1 g178919(.A0 (\cpuregs[5] [28]), .A1 (n_2492), .B0
       (\cpuregs[14] [28]), .B1 (n_2531), .Y (n_2669));
  AOI22X1 g178920(.A0 (\cpuregs[4] [28]), .A1 (n_2529), .B0
       (\cpuregs[3] [28]), .B1 (n_2503), .Y (n_2668));
  AO22X1 g178921(.A0 (\cpuregs[2] [28]), .A1 (n_38), .B0
       (decoded_imm[28]), .B1 (n_421), .Y (n_2667));
  AOI22X1 g178922(.A0 (\cpuregs[6] [28]), .A1 (n_2530), .B0
       (\cpuregs[7] [28]), .B1 (n_12), .Y (n_2666));
  AOI22X1 g178923(.A0 (\cpuregs[12] [28]), .A1 (n_2521), .B0
       (\cpuregs[13] [28]), .B1 (n_2498), .Y (n_2665));
  AOI22X1 g178924(.A0 (\cpuregs[10] [28]), .A1 (n_2520), .B0
       (\cpuregs[11] [28]), .B1 (n_2497), .Y (n_2664));
  AOI22X1 g178925(.A0 (\cpuregs[8] [28]), .A1 (n_2494), .B0
       (\cpuregs[9] [28]), .B1 (n_2526), .Y (n_2663));
  AOI22X1 g178926(.A0 (\cpuregs[29] [28]), .A1 (n_2524), .B0
       (\cpuregs[30] [28]), .B1 (n_2523), .Y (n_2662));
  AOI22X1 g178927(.A0 (\cpuregs[24] [28]), .A1 (n_2490), .B0
       (\cpuregs[23] [28]), .B1 (n_2500), .Y (n_2661));
  AOI22X1 g178928(.A0 (\cpuregs[28] [28]), .A1 (n_2491), .B0
       (\cpuregs[27] [28]), .B1 (n_2525), .Y (n_2660));
  AOI22X1 g178929(.A0 (\cpuregs[25] [28]), .A1 (n_2528), .B0
       (\cpuregs[26] [28]), .B1 (n_2493), .Y (n_2659));
  AOI22X1 g178930(.A0 (\cpuregs[21] [28]), .A1 (n_2495), .B0
       (\cpuregs[22] [28]), .B1 (n_2518), .Y (n_2658));
  AOI22X1 g178931(.A0 (\cpuregs[16] [28]), .A1 (n_2502), .B0
       (\cpuregs[15] [28]), .B1 (n_2504), .Y (n_2657));
  AOI22X1 g178932(.A0 (\cpuregs[20] [28]), .A1 (n_2522), .B0
       (\cpuregs[19] [28]), .B1 (n_2496), .Y (n_2656));
  AOI22X1 g178933(.A0 (\cpuregs[24] [29]), .A1 (n_2490), .B0
       (\cpuregs[23] [29]), .B1 (n_2500), .Y (n_2655));
  AOI22X1 g178934(.A0 (\cpuregs[25] [29]), .A1 (n_2528), .B0
       (\cpuregs[26] [29]), .B1 (n_2493), .Y (n_2654));
  AOI22X1 g178935(.A0 (\cpuregs[29] [29]), .A1 (n_2524), .B0
       (\cpuregs[30] [29]), .B1 (n_2523), .Y (n_2653));
  AOI22X1 g178936(.A0 (\cpuregs[2] [29]), .A1 (n_38), .B0
       (\cpuregs[31] [29]), .B1 (n_2499), .Y (n_2652));
  AOI22X1 g178937(.A0 (\cpuregs[4] [29]), .A1 (n_2529), .B0
       (\cpuregs[5] [29]), .B1 (n_2492), .Y (n_2651));
  AOI22X1 g178938(.A0 (\cpuregs[20] [29]), .A1 (n_2522), .B0
       (\cpuregs[19] [29]), .B1 (n_2496), .Y (n_2650));
  AOI22X1 g178939(.A0 (\cpuregs[16] [29]), .A1 (n_2502), .B0
       (\cpuregs[15] [29]), .B1 (n_2504), .Y (n_2649));
  AOI22X1 g178940(.A0 (\cpuregs[17] [29]), .A1 (n_2527), .B0
       (\cpuregs[18] [29]), .B1 (n_2519), .Y (n_2648));
  AO22X1 g178941(.A0 (\cpuregs[10] [29]), .A1 (n_2520), .B0
       (\cpuregs[7] [29]), .B1 (n_12), .Y (n_2647));
  AOI22X1 g178942(.A0 (\cpuregs[6] [29]), .A1 (n_2530), .B0
       (\reg_op2[29]_9698 ), .B1 (n_832), .Y (n_2646));
  AOI22X1 g178943(.A0 (\cpuregs[12] [29]), .A1 (n_2521), .B0
       (\cpuregs[13] [29]), .B1 (n_2498), .Y (n_2645));
  AOI22X1 g178944(.A0 (\cpuregs[4] [30]), .A1 (n_2529), .B0
       (\cpuregs[5] [30]), .B1 (n_2492), .Y (n_2644));
  AOI22X1 g178945(.A0 (\cpuregs[2] [30]), .A1 (n_38), .B0
       (\cpuregs[3] [30]), .B1 (n_2503), .Y (n_2643));
  AOI22X1 g178946(.A0 (\cpuregs[11] [30]), .A1 (n_2497), .B0
       (\cpuregs[7] [30]), .B1 (n_12), .Y (n_2642));
  AOI22X1 g178947(.A0 (\cpuregs[10] [30]), .A1 (n_2520), .B0
       (\cpuregs[6] [30]), .B1 (n_2530), .Y (n_2641));
  AOI22X1 g178948(.A0 (\cpuregs[12] [30]), .A1 (n_2521), .B0
       (\cpuregs[13] [30]), .B1 (n_2498), .Y (n_2640));
  AOI22X1 g178949(.A0 (\cpuregs[8] [30]), .A1 (n_2494), .B0
       (\cpuregs[9] [30]), .B1 (n_2526), .Y (n_2639));
  AOI22X1 g178950(.A0 (\cpuregs[28] [17]), .A1 (n_2491), .B0
       (\cpuregs[27] [17]), .B1 (n_2525), .Y (n_2638));
  AOI22X1 g178951(.A0 (\cpuregs[20] [30]), .A1 (n_2522), .B0
       (\cpuregs[21] [30]), .B1 (n_2495), .Y (n_2637));
  AOI22X1 g178952(.A0 (\cpuregs[18] [30]), .A1 (n_2519), .B0
       (\cpuregs[19] [30]), .B1 (n_2496), .Y (n_2636));
  AOI22X1 g178953(.A0 (\cpuregs[22] [30]), .A1 (n_2518), .B0
       (\cpuregs[15] [30]), .B1 (n_2504), .Y (n_2635));
  AOI22X1 g178954(.A0 (\cpuregs[29] [30]), .A1 (n_2524), .B0
       (\cpuregs[30] [30]), .B1 (n_2523), .Y (n_2634));
  AOI22X1 g178955(.A0 (\cpuregs[25] [30]), .A1 (n_2528), .B0
       (\cpuregs[26] [30]), .B1 (n_2493), .Y (n_2633));
  AOI22X1 g178956(.A0 (\cpuregs[28] [30]), .A1 (n_2491), .B0
       (\cpuregs[23] [30]), .B1 (n_2500), .Y (n_2632));
  AOI22X1 g178957(.A0 (\cpuregs[24] [30]), .A1 (n_2490), .B0
       (\cpuregs[27] [30]), .B1 (n_2525), .Y (n_2631));
  AOI22X1 g178958(.A0 (\cpuregs[29] [23]), .A1 (n_2524), .B0
       (\cpuregs[30] [23]), .B1 (n_2523), .Y (n_2630));
  AOI22X1 g178959(.A0 (\cpuregs[4] [31]), .A1 (n_2529), .B0
       (\cpuregs[5] [31]), .B1 (n_2492), .Y (n_2629));
  AOI22X1 g178960(.A0 (\cpuregs[2] [31]), .A1 (n_38), .B0
       (\cpuregs[3] [31]), .B1 (n_2503), .Y (n_2628));
  AOI22X1 g178961(.A0 (\cpuregs[12] [31]), .A1 (n_2521), .B0
       (\cpuregs[6] [31]), .B1 (n_2530), .Y (n_2627));
  AOI22X1 g178962(.A0 (\cpuregs[10] [31]), .A1 (n_2520), .B0
       (\cpuregs[11] [31]), .B1 (n_2497), .Y (n_2626));
  AOI22X1 g178963(.A0 (\cpuregs[8] [31]), .A1 (n_2494), .B0
       (\cpuregs[9] [31]), .B1 (n_2526), .Y (n_2625));
  AOI22X1 g178964(.A0 (\cpuregs[26] [31]), .A1 (n_2493), .B0
       (\cpuregs[30] [31]), .B1 (n_2523), .Y (n_2624));
  AOI22X1 g178965(.A0 (\cpuregs[25] [31]), .A1 (n_2528), .B0
       (\cpuregs[27] [31]), .B1 (n_2525), .Y (n_2623));
  AOI22X1 g178966(.A0 (\cpuregs[29] [31]), .A1 (n_2524), .B0
       (\cpuregs[23] [31]), .B1 (n_2500), .Y (n_2622));
  AOI22X1 g178967(.A0 (\cpuregs[21] [31]), .A1 (n_2495), .B0
       (\cpuregs[22] [31]), .B1 (n_2518), .Y (n_2621));
  AOI22X1 g178968(.A0 (\cpuregs[20] [31]), .A1 (n_2522), .B0
       (\cpuregs[19] [31]), .B1 (n_2496), .Y (n_2620));
  AOI22X1 g178969(.A0 (\cpuregs[16] [31]), .A1 (n_2502), .B0
       (\cpuregs[15] [31]), .B1 (n_2504), .Y (n_2619));
  AOI22X1 g178970(.A0 (\cpuregs[17] [31]), .A1 (n_2527), .B0
       (\cpuregs[18] [31]), .B1 (n_2519), .Y (n_2618));
  AOI22X1 g178971(.A0 (\cpuregs[12] [6]), .A1 (n_2521), .B0
       (\cpuregs[13] [6]), .B1 (n_2498), .Y (n_2617));
  AOI22X1 g178972(.A0 (\cpuregs[6] [6]), .A1 (n_2530), .B0
       (\cpuregs[7] [6]), .B1 (n_12), .Y (n_2616));
  NOR4BX1 g178973(.AN (n_2332), .B (n_317), .C (n_2444), .D (n_2446),
       .Y (n_2615));
  OR4X1 g178974(.A (n_679), .B (n_2320), .C (n_2446), .D (n_953), .Y
       (n_2614));
  OAI222X1 g178975(.A0 (n_595), .A1 (n_828), .B0 (n_548), .B1 (n_2508),
       .C0 (n_615), .C1 (n_792), .Y (n_2613));
  NOR4X1 g178976(.A (n_679), .B (n_2320), .C (n_2447), .D (n_953), .Y
       (n_2612));
  AOI32X1 g178977(.A0 (n_854), .A1 (n_2346), .A2 (n_1951), .B0 (n_627),
       .B1 (n_564), .Y (n_2611));
  OAI211X1 g178978(.A0 (n_2330), .A1 (n_2434), .B0 (n_2323), .C0
       (n_2322), .Y (n_2610));
  NAND4XL g178979(.A (n_437), .B (n_504), .C (n_2445), .D (n_673), .Y
       (n_2609));
  AOI32X1 g178980(.A0 (n_692), .A1 (n_2438), .A2 (n_2434), .B0 (n_317),
       .B1 (n_2439), .Y (n_2822));
  INVX1 g178982(.A (n_2603), .Y (n_2604));
  NAND4XL g178985(.A (mem_rdata_q[5]), .B (mem_rdata_q[4]), .C
       (mem_rdata_q[0]), .D (n_2290), .Y (n_2597));
  OAI2BB1X1 g178987(.A0N (n_6533), .A1N (n_2393), .B0 (n_6559), .Y
       (n_2595));
  AND2X1 g178999(.A (n_552), .B (\cpuregs[1] [6]), .Y (n_2594));
  AND2X1 g179000(.A (n_552), .B (\cpuregs[1] [5]), .Y (n_2593));
  AND2X1 g179009(.A (n_552), .B (\cpuregs[1] [23]), .Y (n_2592));
  AND2X1 g179012(.A (n_552), .B (\cpuregs[1] [17]), .Y (n_2591));
  AND2X1 g179014(.A (n_552), .B (\cpuregs[1] [26]), .Y (n_2590));
  NOR2X1 g179015(.A (n_222), .B (n_2485), .Y (n_2589));
  AND2X1 g179016(.A (n_552), .B (\cpuregs[1] [28]), .Y (n_2588));
  AND2X1 g179017(.A (n_552), .B (\cpuregs[1] [10]), .Y (n_2587));
  NOR2X1 g179020(.A (n_504), .B (n_302), .Y (n_2608));
  NOR4X1 g179021(.A (n_326), .B (n_503), .C (n_440), .D (n_2309), .Y
       (n_2607));
  NAND2X1 g179022(.A (n_2506), .B (n_1589), .Y (n_2606));
  NAND2BX1 g179024(.AN (n_2532), .B (n_2336), .Y (n_2605));
  NAND2X1 g179027(.A (n_2513), .B (n_2437), .Y (n_2603));
  OR2X1 g179029(.A (n_325), .B (n_2532), .Y (n_2602));
  NAND2X1 g179030(.A (latched_rd[0]), .B (n_318), .Y (n_2601));
  NAND2X1 g179031(.A (n_681), .B (n_2482), .Y (n_2600));
  OR2X1 g179032(.A (n_2317), .B (n_2506), .Y (n_2599));
  NAND2BX1 g179033(.AN (latched_rd[0]), .B (n_318), .Y (n_2598));
  NAND3BXL g179034(.AN (n_2164), .B (n_1777), .C (n_2382), .Y (n_2582));
  NAND3BXL g179035(.AN (n_2164), .B (n_1771), .C (n_2381), .Y (n_2581));
  NAND3BXL g179036(.AN (n_2164), .B (n_1772), .C (n_2380), .Y (n_2580));
  NAND3BXL g179037(.AN (n_2164), .B (n_1779), .C (n_2379), .Y (n_2579));
  NAND3BXL g179038(.AN (n_2164), .B (n_1780), .C (n_2378), .Y (n_2578));
  NAND3BXL g179039(.AN (n_2164), .B (n_1783), .C (n_2377), .Y (n_2577));
  AOI221X1 g179040(.A0 (\cpuregs[30] [2]), .A1 (n_1622), .B0
       (\cpuregs[31] [2]), .B1 (n_1592), .C0 (n_2472), .Y (n_2576));
  AOI221X1 g179041(.A0 (\cpuregs[22] [3]), .A1 (n_1603), .B0
       (\cpuregs[23] [3]), .B1 (n_1627), .C0 (n_2471), .Y (n_2575));
  AOI221X1 g179042(.A0 (\cpuregs[30] [4]), .A1 (n_1622), .B0
       (\cpuregs[31] [4]), .B1 (n_1592), .C0 (n_2473), .Y (n_2574));
  OAI2BB1X1 g179043(.A0N (instr_srli), .A1N (n_537), .B0 (n_2481), .Y
       (n_2573));
  OAI21X1 g179044(.A0 (n_690), .A1 (n_2336), .B0 (n_2433), .Y (n_2572));
  NOR4X1 g179045(.A (\reg_op2[12]_9681 ), .B (\reg_op2[11]_9680 ), .C
       (\reg_op2[4]_9673 ), .D (n_2182), .Y (n_2571));
  OAI2BB1X1 g179046(.A0N (instr_slli), .A1N (n_537), .B0 (n_2480), .Y
       (n_2570));
  OAI21X1 g179047(.A0 (n_974), .A1 (n_2435), .B0 (n_2324), .Y (n_2569));
  OAI2BB1X1 g179048(.A0N (n_503), .A1N (n_681), .B0 (n_15), .Y
       (n_2568));
  NOR4X1 g179049(.A (n_1353), .B (n_1347), .C (n_1198), .D (n_2278), .Y
       (n_2567));
  AOI32X1 g179050(.A0 (n_538), .A1 (n_1338), .A2 (n_2315), .B0
       (instr_and), .B1 (n_537), .Y (n_2566));
  AOI32X1 g179051(.A0 (n_538), .A1 (n_1344), .A2 (n_2315), .B0
       (instr_or), .B1 (n_537), .Y (n_2565));
  AOI32X1 g179052(.A0 (n_538), .A1 (n_1337), .A2 (n_2315), .B0
       (instr_xor), .B1 (n_537), .Y (n_2564));
  NAND3BXL g179053(.AN (n_2447), .B (n_2445), .C (n_667), .Y (n_2563));
  AOI32X1 g179054(.A0 (n_538), .A1 (n_1326), .A2 (n_2315), .B0
       (instr_slt), .B1 (n_537), .Y (n_2562));
  AOI32X1 g179055(.A0 (is_alu_reg_reg), .A1 (n_538), .A2 (n_2328), .B0
       (instr_sra), .B1 (n_537), .Y (n_2561));
  OAI32X1 g179056(.A0 (n_622), .A1 (n_537), .A2 (n_2329), .B0 (n_766),
       .B1 (n_538), .Y (n_2560));
  NAND3BXL g179057(.AN (n_2164), .B (n_1770), .C (n_2385), .Y (n_2559));
  AOI221X1 g179058(.A0 (\cpuregs[5] [3]), .A1 (n_1611), .B0
       (\cpuregs[15] [3]), .B1 (n_1593), .C0 (n_2348), .Y (n_2558));
  AOI221X1 g179059(.A0 (\cpuregs[5] [0]), .A1 (n_1611), .B0
       (\cpuregs[15] [0]), .B1 (n_1593), .C0 (n_2351), .Y (n_2557));
  AOI221X1 g179060(.A0 (\cpuregs[5] [1]), .A1 (n_1611), .B0
       (\cpuregs[15] [1]), .B1 (n_1593), .C0 (n_2350), .Y (n_2556));
  AOI221X1 g179061(.A0 (\cpuregs[5] [2]), .A1 (n_1611), .B0
       (\cpuregs[15] [2]), .B1 (n_1593), .C0 (n_2349), .Y (n_2555));
  AOI32X1 g179062(.A0 (n_538), .A1 (n_1323), .A2 (n_2315), .B0
       (instr_add), .B1 (n_537), .Y (n_2554));
  AOI32X1 g179063(.A0 (n_538), .A1 (n_1321), .A2 (n_2315), .B0
       (instr_sll), .B1 (n_537), .Y (n_2553));
  AOI32X1 g179064(.A0 (n_538), .A1 (n_1325), .A2 (n_2315), .B0
       (instr_srl), .B1 (n_537), .Y (n_2552));
  MX2X1 g179065(.A (mem_rdata[16]), .B (mem_16bit_buffer[0]), .S0
       (n_431), .Y (n_2551));
  MX2X1 g179066(.A (mem_rdata[17]), .B (mem_16bit_buffer[1]), .S0
       (n_431), .Y (n_2550));
  MX2X1 g179067(.A (mem_rdata[18]), .B (mem_16bit_buffer[2]), .S0
       (n_431), .Y (n_2549));
  MX2X1 g179068(.A (mem_rdata[19]), .B (mem_16bit_buffer[3]), .S0
       (n_431), .Y (n_2548));
  MX2X1 g179069(.A (mem_rdata[20]), .B (mem_16bit_buffer[4]), .S0
       (n_431), .Y (n_2547));
  MX2X1 g179070(.A (mem_rdata[21]), .B (mem_16bit_buffer[5]), .S0
       (n_431), .Y (n_2546));
  MX2X1 g179071(.A (mem_rdata[22]), .B (mem_16bit_buffer[6]), .S0
       (n_431), .Y (n_2545));
  MX2X1 g179072(.A (mem_rdata[23]), .B (mem_16bit_buffer[7]), .S0
       (n_431), .Y (n_2544));
  MX2X1 g179073(.A (mem_rdata[24]), .B (mem_16bit_buffer[8]), .S0
       (n_431), .Y (n_2543));
  MX2X1 g179074(.A (mem_rdata[25]), .B (mem_16bit_buffer[9]), .S0
       (n_431), .Y (n_2542));
  MX2X1 g179075(.A (mem_rdata[26]), .B (mem_16bit_buffer[10]), .S0
       (n_431), .Y (n_2541));
  MX2X1 g179076(.A (mem_rdata[27]), .B (mem_16bit_buffer[11]), .S0
       (n_431), .Y (n_2540));
  MX2X1 g179077(.A (mem_rdata[28]), .B (mem_16bit_buffer[12]), .S0
       (n_431), .Y (n_2539));
  MX2X1 g179078(.A (mem_rdata[29]), .B (mem_16bit_buffer[13]), .S0
       (n_431), .Y (n_2538));
  MX2X1 g179079(.A (mem_rdata[30]), .B (mem_16bit_buffer[14]), .S0
       (n_431), .Y (n_2537));
  MX2X1 g179080(.A (mem_rdata[31]), .B (mem_16bit_buffer[15]), .S0
       (n_431), .Y (n_2536));
  NOR4BX1 g179081(.AN (n_973), .B (is_slli_srli_srai), .C
       (is_jalr_addi_slti_sltiu_xori_ori_andi), .D (n_2327), .Y
       (n_2586));
  NAND2BX1 g179082(.AN (n_14), .B (n_2510), .Y (n_2585));
  NAND3X1 g179083(.A (n_2131), .B (n_2439), .C (n_1619), .Y (n_2584));
  NOR4X1 g179084(.A (n_504), .B (n_334), .C (n_437), .D (n_2320), .Y
       (n_429));
  INVX1 g179085(.A (n_2533), .Y (n_2534));
  NOR2X1 g179086(.A (n_2333), .B (n_325), .Y (n_2517));
  OR4X1 g179088(.A (\genblk2.pcpi_div_quotient_msk [13]), .B
       (\genblk2.pcpi_div_quotient_msk [12]), .C
       (\genblk2.pcpi_div_quotient_msk [11]), .D (n_2157), .Y (n_2516));
  NAND2X1 g179089(.A (n_2316), .B (n_2423), .Y (n_2515));
  NAND2X1 g179090(.A (n_440), .B (n_325), .Y (n_2514));
  NAND2X1 g179092(.A (n_317), .B (n_2436), .Y (n_2535));
  NAND2X1 g179094(.A (n_2439), .B (n_419), .Y (n_2533));
  NAND2X1 g179116(.A (n_2433), .B (n_1588), .Y (n_2532));
  AND2X1 g179138(.A (n_1597), .B (n_344), .Y (n_2531));
  NOR2X4 g179139(.A (n_1623), .B (n_691), .Y (n_2530));
  NOR2X4 g179140(.A (n_1617), .B (n_691), .Y (n_2529));
  AND2X2 g179142(.A (n_1594), .B (n_344), .Y (n_2528));
  AND2X2 g179143(.A (n_1625), .B (n_344), .Y (n_2527));
  AND2X2 g179144(.A (n_1591), .B (n_344), .Y (n_2526));
  AND2X2 g179145(.A (n_1598), .B (n_344), .Y (n_2525));
  AND2X2 g179146(.A (n_1599), .B (n_344), .Y (n_2524));
  AND2X2 g179147(.A (n_1622), .B (n_344), .Y (n_2523));
  NOR2X4 g179148(.A (n_1615), .B (n_691), .Y (n_2522));
  NOR2X4 g179149(.A (n_1609), .B (n_691), .Y (n_2521));
  NOR2X4 g179150(.A (n_1600), .B (n_691), .Y (n_2520));
  AND2X2 g179151(.A (n_10), .B (n_344), .Y (n_2519));
  AND2X2 g179152(.A (n_1603), .B (n_344), .Y (n_2518));
  INVX1 g179155(.A (n_17), .Y (n_2505));
  NAND3X1 g179157(.A (n_1787), .B (n_37), .C (n_2218), .Y (n_2488));
  MX2X1 g179158(.A (mem_wordsize[1]), .B (n_1558), .S0 (n_2325), .Y
       (n_2487));
  MX2X1 g179159(.A (mem_wordsize[0]), .B (n_1557), .S0 (n_2325), .Y
       (n_2486));
  AOI33XL g179160(.A0 (n_582), .A1 (n_901), .A2 (n_2152), .B0 (n_654),
       .B1 (prefetched_high_word), .B2 (n_1862), .Y (n_2485));
  AOI22X1 g179161(.A0 (cpu_state[5]), .A1 (n_2189), .B0 (cpu_state[3]),
       .B1 (n_219), .Y (n_2484));
  NAND4XL g179162(.A (is_alu_reg_reg), .B (n_538), .C (n_1323), .D
       (n_2153), .Y (n_2483));
  NOR4X1 g179163(.A (n_2146), .B (n_2144), .C (n_326), .D (n_503), .Y
       (n_2482));
  NAND4XL g179164(.A (is_alu_reg_imm), .B (n_538), .C (n_1325), .D
       (n_323), .Y (n_2481));
  NAND4XL g179165(.A (is_alu_reg_imm), .B (n_538), .C (n_1321), .D
       (n_323), .Y (n_2480));
  NAND4XL g179166(.A (mem_rdata_q[15]), .B (n_586), .C (n_1321), .D
       (n_1976), .Y (n_2479));
  OAI211X1 g179167(.A0 (n_774), .A1 (n_667), .B0 (n_2335), .C0 (n_355),
       .Y (n_2478));
  OAI211X1 g179168(.A0 (n_685), .A1 (n_342), .B0 (n_1280), .C0 (n_355),
       .Y (n_2477));
  OAI211X1 g179169(.A0 (n_686), .A1 (n_335), .B0 (n_1266), .C0
       (n_2174), .Y (n_2476));
  OAI211X1 g179170(.A0 (n_688), .A1 (n_342), .B0 (n_1233), .C0 (n_355),
       .Y (n_2475));
  OAI221X1 g179171(.A0 (n_564), .A1 (n_1411), .B0 (n_565), .B1 (n_611),
       .C0 (n_2390), .Y (n_2474));
  NAND4XL g179172(.A (n_1869), .B (n_2012), .C (n_2072), .D (n_2306),
       .Y (n_2473));
  NAND4XL g179173(.A (n_1863), .B (n_2062), .C (n_2027), .D (n_2308),
       .Y (n_2472));
  NAND4XL g179174(.A (n_1866), .B (n_2020), .C (n_2021), .D (n_2307),
       .Y (n_2471));
  OAI2BB1X1 g179175(.A0N (n_2319), .A1N (n_1620), .B0 (n_276), .Y
       (n_2470));
  NAND3BXL g179176(.AN (n_2164), .B (n_1774), .C (n_2222), .Y (n_2469));
  NAND3X1 g179177(.A (n_1713), .B (n_1446), .C (n_2192), .Y (n_2468));
  NAND3X1 g179178(.A (n_1454), .B (n_1797), .C (n_2193), .Y (n_2467));
  NAND3X1 g179179(.A (n_1438), .B (n_1939), .C (n_2217), .Y (n_2466));
  NAND3X1 g179180(.A (n_37), .B (n_1795), .C (n_2272), .Y (n_2465));
  NAND3X1 g179181(.A (n_37), .B (n_1781), .C (n_2271), .Y (n_2464));
  NAND3X1 g179182(.A (n_37), .B (n_1785), .C (n_2270), .Y (n_2463));
  NAND3X1 g179183(.A (n_37), .B (n_1789), .C (n_2269), .Y (n_2462));
  NAND3X1 g179184(.A (n_37), .B (n_1791), .C (n_2268), .Y (n_2461));
  NAND3X1 g179185(.A (n_37), .B (n_1793), .C (n_2267), .Y (n_2460));
  NAND3X1 g179186(.A (n_37), .B (n_1792), .C (n_2266), .Y (n_2459));
  NAND3X1 g179187(.A (n_37), .B (n_1794), .C (n_2265), .Y (n_2458));
  NAND3X1 g179188(.A (n_37), .B (n_1768), .C (n_2264), .Y (n_2457));
  NAND3X1 g179189(.A (n_37), .B (n_1790), .C (n_2263), .Y (n_2456));
  NAND3X1 g179190(.A (n_37), .B (n_1786), .C (n_2221), .Y (n_2455));
  NAND3X1 g179191(.A (n_1447), .B (n_1800), .C (n_2194), .Y (n_2454));
  NAND3X1 g179192(.A (n_37), .B (n_1788), .C (n_2220), .Y (n_2453));
  NAND3X1 g179193(.A (n_37), .B (n_1756), .C (n_2219), .Y (n_2452));
  NAND3X1 g179194(.A (n_37), .B (n_1784), .C (n_2260), .Y (n_2451));
  NAND3X1 g179195(.A (n_1456), .B (n_1938), .C (n_2195), .Y (n_2450));
  NAND2X1 g179196(.A (n_2435), .B (n_1620), .Y (n_2513));
  NOR4X1 g179199(.A (cpu_state[6]), .B (n_852), .C (cpu_state[3]), .D
       (n_11749), .Y (n_2512));
  AOI21X1 g179200(.A0 (n_2318), .A1 (n_419), .B0 (n_2449), .Y (n_2511));
  NAND2X1 g179201(.A (n_2435), .B (n_1330), .Y (n_2510));
  OAI21X1 g179202(.A0 (n_323), .A1 (n_2328), .B0 (n_1634), .Y (n_2509));
  OAI31X1 g179203(.A0 (is_sll_srl_sra), .A1 (is_sb_sh_sw), .A2 (n_305),
       .B0 (n_981), .Y (n_2508));
  NOR4BX1 g179204(.AN (n_11), .B (n_14409_BAR), .C (n_1977), .D
       (n_324), .Y (n_318));
  NOR2X1 g179205(.A (n_11741), .B (n_2434), .Y (n_2506));
  AND2X2 g179209(.A (n_1593), .B (n_344), .Y (n_2504));
  AND2X2 g179210(.A (n_1607), .B (n_344), .Y (n_2503));
  AND2X2 g179211(.A (n_1596), .B (n_344), .Y (n_2502));
  AND2X1 g179212(.A (n_344), .B (n_1626), .Y (n_552));
  AND2X2 g179213(.A (n_1627), .B (n_344), .Y (n_2500));
  AND2X2 g179214(.A (n_1592), .B (n_344), .Y (n_2499));
  AND2X2 g179215(.A (n_1606), .B (n_344), .Y (n_2498));
  AND2X2 g179216(.A (n_1608), .B (n_344), .Y (n_2497));
  AND2X2 g179217(.A (n_1605), .B (n_344), .Y (n_2496));
  AND2X2 g179218(.A (n_1614), .B (n_344), .Y (n_2495));
  AND2X2 g179219(.A (n_1595), .B (n_344), .Y (n_2494));
  NOR2X4 g179220(.A (n_11745), .B (n_691), .Y (n_2493));
  AND2X2 g179221(.A (n_1611), .B (n_344), .Y (n_2492));
  AND2X2 g179222(.A (n_9), .B (n_344), .Y (n_2491));
  AND2X2 g179223(.A (n_1604), .B (n_344), .Y (n_2490));
  OR2X1 g179224(.A (n_659), .B (n_2391), .Y (n_2489));
  INVX1 g179225(.A (n_2448), .Y (n_2449));
  INVX1 g179226(.A (n_2444), .Y (n_2445));
  INVX1 g179227(.A (n_2442), .Y (n_2441));
  INVX1 g179229(.A (n_2439), .Y (n_2438));
  INVX1 g179230(.A (n_2437), .Y (n_2436));
  INVX1 g179232(.A (n_2434), .Y (n_2433));
  NOR2X1 g179234(.A (n_544), .B (n_2186), .Y (n_2431));
  NOR2BX1 g179235(.AN (n_2326), .B (mem_do_rinst), .Y (n_2430));
  NOR2X1 g179236(.A (n_544), .B (n_2184), .Y (n_2429));
  NOR2X1 g179237(.A (n_544), .B (n_2185), .Y (n_2428));
  NOR2X1 g179238(.A (n_853), .B (n_2314), .Y (n_2427));
  NAND2X1 g179269(.A (n_2324), .B (n_1588), .Y (n_2448));
  NAND2X1 g179274(.A (n_680), .B (n_2337), .Y (n_2447));
  NAND2X1 g179276(.A (n_504), .B (n_2337), .Y (n_2446));
  NAND2X1 g179307(.A (n_679), .B (n_2333), .Y (n_2444));
  NAND2X1 g179310(.A (n_2317), .B (n_419), .Y (n_2443));
  NAND2X1 g179311(.A (cpu_state[5]), .B (n_2327), .Y (n_2442));
  NOR2X1 g179313(.A (n_685), .B (n_2316), .Y (n_2440));
  NOR2X1 g179314(.A (n_438), .B (n_2316), .Y (n_2439));
  NAND2X1 g179315(.A (n_2324), .B (n_1589), .Y (n_2437));
  NOR2X1 g179316(.A (n_687), .B (n_2319), .Y (n_2435));
  NAND2X1 g179317(.A (n_327), .B (n_2332), .Y (n_2434));
  AND2X2 g179318(.A (n_659), .B (n_2327), .Y (n_344));
  INVX1 g179319(.A (n_2425), .Y (n_2426));
  INVX1 g179320(.A (n_2422), .Y (n_2421));
  MX2X1 g179322(.A (n_1953), .B (mem_do_rdata), .S0 (n_2155), .Y
       (n_2418));
  OAI222X1 g179323(.A0 (n_680), .A1 (n_335), .B0 (n_1804), .B1 (n_342),
       .C0 (n_733), .C1 (n_667), .Y (n_2417));
  OAI222X1 g179324(.A0 (n_683), .A1 (n_335), .B0 (n_1808), .B1 (n_342),
       .C0 (n_772), .C1 (n_667), .Y (n_2416));
  AOI2BB1X1 g179325(.A0N (n_767), .A1N (n_305), .B0
       (is_slli_srli_srai), .Y (n_2415));
  NAND4XL g179326(.A (mem_valid_9465), .B (n_1341), .C (n_1956), .D
       (n_1918), .Y (n_2414));
  OAI211X1 g179328(.A0 (n_731), .A1 (n_667), .B0 (n_2168), .C0 (n_355),
       .Y (n_2412));
  OAI211X1 g179329(.A0 (n_775), .A1 (n_667), .B0 (n_2167), .C0 (n_355),
       .Y (n_2411));
  OAI211X1 g179330(.A0 (n_588), .A1 (n_540), .B0 (n_903), .C0 (n_36),
       .Y (n_2410));
  OAI211X1 g179331(.A0 (n_590), .A1 (n_540), .B0 (n_949), .C0 (n_36),
       .Y (n_2409));
  OAI211X1 g179332(.A0 (n_648), .A1 (n_540), .B0 (n_936), .C0 (n_36),
       .Y (n_2408));
  OAI211X1 g179333(.A0 (n_591), .A1 (n_540), .B0 (n_805), .C0 (n_36),
       .Y (n_2407));
  OAI211X1 g179334(.A0 (n_727), .A1 (n_540), .B0 (n_906), .C0 (n_36),
       .Y (n_2406));
  OAI211X1 g179335(.A0 (n_752), .A1 (n_540), .B0 (n_827), .C0 (n_36),
       .Y (n_2405));
  NAND3BXL g179336(.AN (n_2169), .B (n_1278), .C (n_355), .Y (n_2404));
  OAI211X1 g179337(.A0 (n_644), .A1 (n_540), .B0 (n_798), .C0 (n_36),
       .Y (n_2403));
  OAI211X1 g179338(.A0 (n_581), .A1 (n_540), .B0 (n_945), .C0 (n_36),
       .Y (n_2402));
  OAI211X1 g179339(.A0 (n_579), .A1 (n_540), .B0 (n_911), .C0 (n_36),
       .Y (n_2401));
  OAI211X1 g179340(.A0 (n_639), .A1 (n_540), .B0 (n_887), .C0 (n_36),
       .Y (n_2400));
  OAI211X1 g179341(.A0 (n_642), .A1 (n_540), .B0 (n_819), .C0 (n_36),
       .Y (n_2399));
  OAI211X1 g179342(.A0 (n_771), .A1 (n_667), .B0 (n_2173), .C0 (n_355),
       .Y (n_2398));
  OAI222X1 g179343(.A0 (n_689), .A1 (n_335), .B0 (n_1816), .B1 (n_342),
       .C0 (n_769), .C1 (n_667), .Y (n_2397));
  OAI211X1 g179344(.A0 (n_636), .A1 (n_540), .B0 (n_923), .C0 (n_36),
       .Y (n_2396));
  OAI211X1 g179345(.A0 (n_679), .A1 (n_335), .B0 (n_1259), .C0
       (n_2172), .Y (n_2395));
  OAI211X1 g179346(.A0 (n_1809), .A1 (n_342), .B0 (n_1254), .C0
       (n_355), .Y (n_2394));
  OAI211X1 g179347(.A0 (n_629), .A1 (n_1914), .B0 (n_6537), .C0
       (n_7145), .Y (n_2393));
  AOI21X1 g179348(.A0 (reg_sh[3]), .A1 (n_2151), .B0 (n_2338), .Y
       (n_2392));
  OAI31X1 g179349(.A0 (n_611), .A1 (n_1955), .A2 (n_544), .B0 (n_2166),
       .Y (n_2391));
  OAI211X1 g179350(.A0 (cpu_state[5]), .A1 (n_54), .B0 (n_14409_BAR),
       .C0 (n_2128), .Y (n_2390));
  OAI221X1 g179351(.A0 (n_637), .A1 (n_677), .B0 (n_747), .B1 (n_1940),
       .C0 (n_2183), .Y (n_2389));
  OAI2BB1X1 g179352(.A0N (n_14409_BAR), .A1N (n_297), .B0 (n_613), .Y
       (n_2388));
  OAI211X1 g179353(.A0 (n_735), .A1 (n_667), .B0 (n_2176), .C0 (n_355),
       .Y (n_2387));
  AOI222X1 g179354(.A0 (\reg_op1[5]_9642 ), .A1 (n_550), .B0
       (\reg_op1[3]_9640 ), .B1 (n_1941), .C0 (n_833), .C1 (n_6956), .Y
       (n_2386));
  AOI222X1 g179355(.A0 (cpu_state[3]), .A1 (n_72), .B0 (n_1720), .B1
       (cpu_state[5]), .C0 (\reg_op1[9]_9646 ), .C1 (cpu_state[2]), .Y
       (n_2385));
  OAI211X1 g179356(.A0 (n_643), .A1 (n_875), .B0 (n_2124), .C0
       (n_1443), .Y (n_2384));
  OAI222X1 g179357(.A0 (n_2145), .A1 (n_335), .B0 (n_1806), .B1
       (n_342), .C0 (n_776), .C1 (n_667), .Y (n_2383));
  AOI222X1 g179358(.A0 (cpu_state[3]), .A1 (n_70), .B0 (n_1715), .B1
       (cpu_state[5]), .C0 (\reg_op1[8]_9645 ), .C1 (cpu_state[2]), .Y
       (n_2382));
  AOI222X1 g179359(.A0 (cpu_state[3]), .A1 (n_74), .B0 (n_1714), .B1
       (cpu_state[5]), .C0 (\reg_op1[10]_9647 ), .C1 (cpu_state[2]), .Y
       (n_2381));
  AOI222X1 g179360(.A0 (cpu_state[3]), .A1 (n_78), .B0 (n_1727), .B1
       (cpu_state[5]), .C0 (\reg_op1[11]_9648 ), .C1 (cpu_state[2]), .Y
       (n_2380));
  AOI222X1 g179361(.A0 (cpu_state[3]), .A1 (n_76), .B0 (n_1801), .B1
       (cpu_state[5]), .C0 (\reg_op1[12]_9649 ), .C1 (cpu_state[2]), .Y
       (n_2379));
  AOI222X1 g179362(.A0 (cpu_state[3]), .A1 (n_80), .B0 (n_1722), .B1
       (cpu_state[5]), .C0 (\reg_op1[13]_9650 ), .C1 (cpu_state[2]), .Y
       (n_2378));
  AOI222X1 g179363(.A0 (cpu_state[3]), .A1 (n_84), .B0 (n_1712), .B1
       (n_1183), .C0 (\reg_op1[14]_9651 ), .C1 (cpu_state[2]), .Y
       (n_2377));
  OAI211X1 g179368(.A0 (n_681), .A1 (n_335), .B0 (n_1261), .C0
       (n_2170), .Y (n_2372));
  OAI221X1 g179369(.A0 (n_564), .A1 (n_1523), .B0 (n_744), .B1 (n_611),
       .C0 (n_2191), .Y (n_2371));
  AOI222X1 g179370(.A0 (\reg_op1[25]_9662 ), .A1 (n_550), .B0
       (\reg_op1[23]_9660 ), .B1 (n_1941), .C0 (n_833), .C1 (n_6936),
       .Y (n_2370));
  AOI222X1 g179371(.A0 (\reg_op1[27]_9664 ), .A1 (n_550), .B0
       (\reg_op1[25]_9662 ), .B1 (n_1941), .C0 (n_833), .C1 (n_6934),
       .Y (n_2369));
  AOI222X1 g179372(.A0 (\reg_op1[28]_9665 ), .A1 (n_550), .B0
       (\reg_op1[26]_9663 ), .B1 (n_1941), .C0 (n_833), .C1 (n_6933),
       .Y (n_2368));
  AOI222X1 g179373(.A0 (\reg_op1[29]_9666 ), .A1 (n_550), .B0
       (\reg_op1[27]_9664 ), .B1 (n_1941), .C0 (n_833), .C1 (n_6932),
       .Y (n_2367));
  OAI2BB1X1 g179374(.A0N (n_503), .A1N (n_674), .B0 (n_2198), .Y
       (n_2366));
  AOI222X1 g179375(.A0 (\reg_op1[6]_9643 ), .A1 (n_550), .B0
       (\reg_op1[4]_9641 ), .B1 (n_1941), .C0 (n_833), .C1 (n_6955), .Y
       (n_2365));
  AOI222X1 g179376(.A0 (\reg_op1[7]_9644 ), .A1 (n_550), .B0
       (\reg_op1[5]_9642 ), .B1 (n_1941), .C0 (n_833), .C1 (n_6954), .Y
       (n_2364));
  MX2X1 g179377(.A (is_jalr_addi_slti_sltiu_xori_ori_andi), .B
       (n_2126), .S0 (n_538), .Y (n_2363));
  AOI222X1 g179378(.A0 (\reg_op1[16]_9653 ), .A1 (n_550), .B0
       (\reg_op1[14]_9651 ), .B1 (n_1941), .C0 (n_833), .C1 (n_6945),
       .Y (n_2362));
  AOI222X1 g179379(.A0 (\reg_op1[18]_9655 ), .A1 (n_550), .B0
       (\reg_op1[16]_9653 ), .B1 (n_1941), .C0 (n_833), .C1 (n_6943),
       .Y (n_2361));
  AOI222X1 g179380(.A0 (\reg_op1[14]_9651 ), .A1 (n_550), .B0
       (\reg_op1[12]_9649 ), .B1 (n_1941), .C0 (n_833), .C1 (n_6947),
       .Y (n_2360));
  AOI222X1 g179381(.A0 (\reg_op1[12]_9649 ), .A1 (n_550), .B0
       (\reg_op1[10]_9647 ), .B1 (n_1941), .C0 (n_833), .C1 (n_6949),
       .Y (n_2359));
  AOI222X1 g179382(.A0 (\reg_op1[13]_9650 ), .A1 (n_550), .B0
       (\reg_op1[11]_9648 ), .B1 (n_1941), .C0 (n_833), .C1 (n_6948),
       .Y (n_2358));
  AOI222X1 g179383(.A0 (\reg_op1[9]_9646 ), .A1 (n_550), .B0
       (\reg_op1[7]_9644 ), .B1 (n_1941), .C0 (n_833), .C1 (n_6952), .Y
       (n_2357));
  AOI222X1 g179384(.A0 (\reg_op1[10]_9647 ), .A1 (n_550), .B0
       (\reg_op1[8]_9645 ), .B1 (n_1941), .C0 (n_833), .C1 (n_6951), .Y
       (n_2356));
  AOI222X1 g179385(.A0 (\reg_op1[11]_9648 ), .A1 (n_550), .B0
       (\reg_op1[9]_9646 ), .B1 (n_1941), .C0 (n_833), .C1 (n_6950), .Y
       (n_2355));
  OAI21X1 g179386(.A0 (n_2143), .A1 (n_335), .B0 (n_2261), .Y (n_2354));
  NAND4XL g179387(.A (n_2039), .B (n_2038), .C (n_2056), .D (n_2059),
       .Y (n_2353));
  NAND4XL g179388(.A (n_2047), .B (n_2048), .C (n_2046), .D (n_2052),
       .Y (n_2352));
  NAND4XL g179389(.A (n_2042), .B (n_2053), .C (n_2054), .D (n_2043),
       .Y (n_2351));
  NAND4XL g179390(.A (n_2058), .B (n_2035), .C (n_2110), .D (n_2057),
       .Y (n_2350));
  NAND4XL g179391(.A (n_2067), .B (n_2032), .C (n_2030), .D (n_2031),
       .Y (n_2349));
  NAND4XL g179392(.A (n_2025), .B (n_2063), .C (n_2055), .D (n_2024),
       .Y (n_2348));
  NAND4XL g179393(.A (n_2069), .B (n_2017), .C (n_2015), .D (n_2016),
       .Y (n_2347));
  AOI22X1 g179394(.A0 (n_2156), .A1 (mem_rdata[31]), .B0 (n_990), .B1
       (mem_rdata[15]), .Y (n_2346));
  MX2X1 g179395(.A (decoded_imm_j[12]), .B (n_317), .S0 (n_667), .Y
       (n_2345));
  MX2X1 g179396(.A (n_293), .B (mem_do_wdata), .S0 (n_2154), .Y
       (n_2344));
  MX2X1 g179397(.A (mem_rdata_q[2]), .B (n_504), .S0 (n_446), .Y
       (n_2343));
  OAI22X1 g179398(.A0 (n_445), .A1 (n_679), .B0 (n_594), .B1 (n_446),
       .Y (n_2342));
  OAI22X1 g179399(.A0 (n_445), .A1 (n_686), .B0 (n_649), .B1 (n_446),
       .Y (n_2341));
  OAI22X1 g179400(.A0 (n_445), .A1 (n_683), .B0 (n_586), .B1 (n_446),
       .Y (n_2340));
  OAI211X1 g179401(.A0 (n_682), .A1 (n_335), .B0 (n_1269), .C0
       (n_2171), .Y (n_2339));
  NAND2X1 g179402(.A (n_2321), .B (n_1588), .Y (n_2425));
  NAND2X1 g179403(.A (n_2318), .B (n_1620), .Y (n_2424));
  NAND3X1 g179404(.A (n_439), .B (n_438), .C (n_687), .Y (n_2423));
  NAND2X1 g179405(.A (n_2317), .B (n_1620), .Y (n_2422));
  NAND3X1 g179406(.A (n_503), .B (n_440), .C (n_2131), .Y (n_325));
  AND2X1 g179407(.A (n_2293), .B (n_1874), .Y (n_431));
  INVX1 g179409(.A (n_11741), .Y (n_2330));
  INVX1 g179410(.A (n_2328), .Y (n_2329));
  INVX1 g179411(.A (n_2324), .Y (n_2323));
  INVX1 g179412(.A (n_2322), .Y (n_2321));
  INVX1 g179414(.A (n_2319), .Y (n_2318));
  INVX1 g179415(.A (n_2317), .Y (n_2316));
  INVX1 g179416(.A (n_2314), .Y (n_2315));
  AOI21X1 g179418(.A0 (n_787), .A1 (n_1796), .B0 (n_544), .Y (n_2312));
  AOI221X1 g179419(.A0 (\cpuregs[2] [1]), .A1 (n_1621), .B0
       (\cpuregs[23] [1]), .B1 (n_1627), .C0 (n_2040), .Y (n_2311));
  AOI221X1 g179420(.A0 (\cpuregs[1] [0]), .A1 (n_1626), .B0
       (\cpuregs[27] [0]), .B1 (n_1598), .C0 (n_11800), .Y (n_2310));
  NAND2X1 g179421(.A (n_2143), .B (n_2146), .Y (n_2309));
  AOI221X1 g179422(.A0 (\cpuregs[22] [2]), .A1 (n_1603), .B0
       (\cpuregs[23] [2]), .B1 (n_1627), .C0 (n_2028), .Y (n_2308));
  AOI221X1 g179423(.A0 (\cpuregs[28] [3]), .A1 (n_9), .B0
       (\cpuregs[29] [3]), .B1 (n_1599), .C0 (n_2019), .Y (n_2307));
  AOI221X1 g179424(.A0 (\cpuregs[22] [4]), .A1 (n_1603), .B0
       (\cpuregs[23] [4]), .B1 (n_1627), .C0 (n_2011), .Y (n_2306));
  NOR2X1 g179425(.A (n_2009), .B (n_850), .Y (n_2305));
  OAI211X1 g179426(.A0 (n_597), .A1 (n_540), .B0 (n_1425), .C0
       (n_2163), .Y (n_2304));
  OAI211X1 g179427(.A0 (n_596), .A1 (n_540), .B0 (n_1426), .C0
       (n_2163), .Y (n_2303));
  OAI211X1 g179428(.A0 (n_728), .A1 (n_540), .B0 (n_1445), .C0
       (n_2163), .Y (n_2302));
  OAI211X1 g179429(.A0 (n_762), .A1 (n_540), .B0 (n_1427), .C0
       (n_2163), .Y (n_2301));
  OAI211X1 g179430(.A0 (n_583), .A1 (n_540), .B0 (n_1428), .C0
       (n_2163), .Y (n_2300));
  OAI211X1 g179431(.A0 (n_641), .A1 (n_540), .B0 (n_1442), .C0
       (n_2163), .Y (n_2299));
  OAI211X1 g179432(.A0 (n_640), .A1 (n_540), .B0 (n_1455), .C0
       (n_2163), .Y (n_2298));
  NAND2BX1 g179433(.AN (n_1635), .B (n_2127), .Y (n_2297));
  OAI211X1 g179434(.A0 (n_616), .A1 (n_540), .B0 (n_1465), .C0
       (n_2163), .Y (n_2296));
  OAI32X1 g179435(.A0 (n_356), .A1 (n_832), .A2 (n_1535), .B0 (n_793),
       .B1 (n_989), .Y (n_2295));
  NOR2X1 g179436(.A (n_1979), .B (n_544), .Y (n_2294));
  NAND2X1 g179437(.A (n_582), .B (n_2152), .Y (n_2293));
  NOR2X1 g179438(.A (n_1981), .B (n_544), .Y (n_2292));
  NOR2X1 g179439(.A (n_1982), .B (n_544), .Y (n_2291));
  NOR4X1 g179440(.A (mem_rdata_q[18]), .B (mem_rdata_q[19]), .C
       (mem_rdata_q[17]), .D (n_1534), .Y (n_2290));
  NOR2X1 g179441(.A (n_1997), .B (n_544), .Y (n_2289));
  NOR2X1 g179442(.A (n_1985), .B (n_544), .Y (n_2288));
  NOR2X1 g179443(.A (n_1986), .B (n_544), .Y (n_2287));
  NOR2X1 g179444(.A (n_1987), .B (n_544), .Y (n_2286));
  NOR2X1 g179445(.A (n_1989), .B (n_544), .Y (n_2285));
  NOR2X1 g179446(.A (n_1993), .B (n_544), .Y (n_2284));
  NOR2X1 g179447(.A (n_1988), .B (n_544), .Y (n_2283));
  NOR2X1 g179448(.A (n_1994), .B (n_544), .Y (n_2282));
  OAI211X1 g179449(.A0 (n_947), .A1 (n_119), .B0 (n_1915), .C0
       (n_1974), .Y (n_2281));
  OAI211X1 g179456(.A0 (n_278), .A1 (n_1195), .B0 (n_1305), .C0
       (n_1408), .Y (n_2280));
  NOR2X1 g179465(.A (reg_sh[3]), .B (n_2151), .Y (n_2338));
  NOR2X1 g179469(.A (n_276), .B (n_437), .Y (n_2337));
  NOR2X1 g179484(.A (n_317), .B (n_440), .Y (n_2336));
  NAND2X1 g179493(.A (n_327), .B (n_673), .Y (n_2335));
  NAND2BX1 g179495(.AN (n_305), .B (is_sb_sh_sw), .Y (n_2334));
  NOR2X1 g179496(.A (n_683), .B (n_686), .Y (n_2333));
  NOR2X1 g179499(.A (n_439), .B (n_438), .Y (n_2332));
  AND2X1 g179503(.A (n_2153), .B (n_1325), .Y (n_2328));
  NAND2X1 g179505(.A (n_356), .B (n_305), .Y (n_2327));
  OAI211X1 g179506(.A0 (n_6567), .A1 (n_664), .B0 (n_1956), .C0
       (n_1957), .Y (n_2326));
  NAND2X1 g179509(.A (n_324), .B (n_2166), .Y (n_2325));
  NOR2X1 g179510(.A (n_685), .B (n_687), .Y (n_2324));
  NAND2X1 g179513(.A (n_439), .B (n_685), .Y (n_2322));
  NAND2X1 g179514(.A (n_686), .B (n_683), .Y (n_2320));
  NAND2X1 g179515(.A (n_438), .B (n_688), .Y (n_2319));
  NOR2X1 g179516(.A (n_439), .B (n_327), .Y (n_2317));
  NAND2X1 g179517(.A (is_alu_reg_reg), .B (n_323), .Y (n_2314));
  NAND2X1 g179518(.A (n_317), .B (n_674), .Y (n_355));
  OAI221X1 g179521(.A0 (n_278), .A1 (n_1196), .B0 (n_916), .B1 (n_119),
       .C0 (n_1416), .Y (n_2279));
  NAND4XL g179522(.A (n_1194), .B (n_1359), .C (n_1360), .D (n_1559),
       .Y (n_2278));
  OAI211X1 g179523(.A0 (n_590), .A1 (n_34), .B0 (n_1537), .C0 (n_1488),
       .Y (n_2277));
  OAI221X1 g179524(.A0 (n_644), .A1 (n_34), .B0 (n_647), .B1 (n_1327),
       .C0 (n_1464), .Y (n_2276));
  OAI221X1 g179525(.A0 (n_581), .A1 (n_34), .B0 (n_650), .B1 (n_1327),
       .C0 (n_1460), .Y (n_2275));
  OAI211X1 g179526(.A0 (n_639), .A1 (n_34), .B0 (n_1532), .C0 (n_1476),
       .Y (n_2274));
  OAI32X1 g179527(.A0 (n_982), .A1 (n_854), .A2 (n_676), .B0 (n_716),
       .B1 (n_1940), .Y (n_2273));
  AOI22X1 g179528(.A0 (n_1738), .A1 (n_1181), .B0 (\reg_op1[21]_9658 ),
       .B1 (cpu_state[2]), .Y (n_2272));
  AOI22X1 g179529(.A0 (n_1726), .A1 (n_1190), .B0 (\reg_op1[22]_9659 ),
       .B1 (cpu_state[2]), .Y (n_2271));
  AOI22X1 g179530(.A0 (n_1737), .A1 (n_1174), .B0 (\reg_op1[23]_9660 ),
       .B1 (cpu_state[2]), .Y (n_2270));
  AOI22X1 g179531(.A0 (n_1736), .A1 (n_1188), .B0 (\reg_op1[24]_9661 ),
       .B1 (cpu_state[2]), .Y (n_2269));
  AOI22X1 g179532(.A0 (n_1735), .A1 (n_1173), .B0 (\reg_op1[25]_9662 ),
       .B1 (cpu_state[2]), .Y (n_2268));
  AOI22X1 g179533(.A0 (n_1728), .A1 (n_1185), .B0 (\reg_op1[26]_9663 ),
       .B1 (cpu_state[2]), .Y (n_2267));
  AOI22X1 g179534(.A0 (n_1734), .A1 (n_1178), .B0 (\reg_op1[27]_9664 ),
       .B1 (cpu_state[2]), .Y (n_2266));
  AOI22X1 g179535(.A0 (n_1733), .A1 (n_1169), .B0 (\reg_op1[28]_9665 ),
       .B1 (cpu_state[2]), .Y (n_2265));
  AOI22X1 g179536(.A0 (n_1716), .A1 (n_1187), .B0 (\reg_op1[29]_9666 ),
       .B1 (cpu_state[2]), .Y (n_2264));
  AOI22X1 g179537(.A0 (n_1732), .A1 (n_1168), .B0 (\reg_op1[30]_9667 ),
       .B1 (cpu_state[2]), .Y (n_2263));
  OAI2BB1X1 g179538(.A0N (\genblk1.pcpi_mul_rs1 [32]), .A1N (n_672),
       .B0 (n_2123), .Y (n_2262));
  AOI22X1 g179539(.A0 (n_1814), .A1 (n_673), .B0 (decoded_imm_j[8]),
       .B1 (n_953), .Y (n_2261));
  AOI22X1 g179540(.A0 (n_1739), .A1 (n_1170), .B0 (\reg_op1[20]_9657 ),
       .B1 (cpu_state[2]), .Y (n_2260));
  OAI222X1 g179541(.A0 (n_776), .A1 (n_662), .B0 (n_579), .B1 (n_1947),
       .C0 (n_732), .C1 (n_538), .Y (n_2259));
  OAI2BB1X1 g179542(.A0N (mem_rdata_q[29]), .A1N (n_1946), .B0
       (n_1433), .Y (n_2258));
  OAI2BB1X1 g179543(.A0N (n_6574), .A1N (n_353), .B0 (n_2103), .Y
       (n_2257));
  OAI2BB1X1 g179544(.A0N (n_6575), .A1N (n_353), .B0 (n_2102), .Y
       (n_2256));
  OAI2BB1X1 g179545(.A0N (n_6576), .A1N (n_353), .B0 (n_2101), .Y
       (n_2255));
  OAI2BB1X1 g179546(.A0N (n_6577), .A1N (n_353), .B0 (n_2100), .Y
       (n_2254));
  OAI2BB1X1 g179547(.A0N (n_6578), .A1N (n_353), .B0 (n_2099), .Y
       (n_2253));
  OAI2BB1X1 g179548(.A0N (n_353), .A1N (n_6579), .B0 (n_2098), .Y
       (n_2252));
  OAI2BB1X1 g179549(.A0N (n_353), .A1N (n_6580), .B0 (n_2097), .Y
       (n_2251));
  OAI2BB1X1 g179550(.A0N (n_353), .A1N (n_6581), .B0 (n_2096), .Y
       (n_2250));
  OAI2BB1X1 g179551(.A0N (n_353), .A1N (n_6582), .B0 (n_2095), .Y
       (n_2249));
  OAI2BB1X1 g179552(.A0N (n_353), .A1N (n_6583), .B0 (n_2094), .Y
       (n_2248));
  OAI2BB1X1 g179553(.A0N (n_353), .A1N (n_6584), .B0 (n_2093), .Y
       (n_2247));
  OAI2BB1X1 g179554(.A0N (n_353), .A1N (n_6585), .B0 (n_2092), .Y
       (n_2246));
  OAI2BB1X1 g179555(.A0N (n_353), .A1N (n_6586), .B0 (n_2091), .Y
       (n_2245));
  OAI2BB1X1 g179556(.A0N (n_353), .A1N (n_6587), .B0 (n_2090), .Y
       (n_2244));
  OAI2BB1X1 g179557(.A0N (n_353), .A1N (n_6588), .B0 (n_2089), .Y
       (n_2243));
  OAI2BB1X1 g179558(.A0N (n_353), .A1N (n_6589), .B0 (n_2088), .Y
       (n_2242));
  OAI2BB1X1 g179559(.A0N (n_353), .A1N (n_6590), .B0 (n_2087), .Y
       (n_2241));
  OAI2BB1X1 g179560(.A0N (n_353), .A1N (n_6591), .B0 (n_2086), .Y
       (n_2240));
  OAI2BB1X1 g179561(.A0N (n_353), .A1N (n_6593), .B0 (n_2084), .Y
       (n_2239));
  OAI2BB1X1 g179562(.A0N (n_353), .A1N (n_6594), .B0 (n_2083), .Y
       (n_2238));
  OAI2BB1X1 g179563(.A0N (n_353), .A1N (n_6595), .B0 (n_2082), .Y
       (n_2237));
  OAI2BB1X1 g179564(.A0N (n_353), .A1N (n_6596), .B0 (n_2081), .Y
       (n_2236));
  OAI2BB1X1 g179565(.A0N (n_353), .A1N (n_6597), .B0 (n_2080), .Y
       (n_2235));
  OAI2BB1X1 g179566(.A0N (n_353), .A1N (n_6598), .B0 (n_2079), .Y
       (n_2234));
  OAI2BB1X1 g179567(.A0N (n_353), .A1N (n_6600), .B0 (n_2077), .Y
       (n_2233));
  OAI2BB1X1 g179568(.A0N (n_353), .A1N (n_6601), .B0 (n_2076), .Y
       (n_2232));
  OAI2BB1X1 g179569(.A0N (n_353), .A1N (n_6602), .B0 (n_2075), .Y
       (n_2231));
  OAI2BB1X1 g179570(.A0N (n_353), .A1N (n_6603), .B0 (n_2074), .Y
       (n_2230));
  OAI2BB1X1 g179571(.A0N (mem_rdata_q[28]), .A1N (n_1946), .B0
       (n_1462), .Y (n_2229));
  OAI222X1 g179572(.A0 (n_733), .A1 (n_662), .B0 (n_648), .B1 (n_1947),
       .C0 (n_768), .C1 (n_538), .Y (n_2228));
  OAI2BB1X1 g179573(.A0N (n_353), .A1N (n_6604), .B0 (n_2073), .Y
       (n_2227));
  OAI2BB1X1 g179574(.A0N (n_353), .A1N (n_6599), .B0 (n_2078), .Y
       (n_2226));
  OAI2BB1X1 g179575(.A0N (n_353), .A1N (n_6592), .B0 (n_2085), .Y
       (n_2225));
  OAI222X1 g179576(.A0 (n_769), .A1 (n_662), .B0 (n_591), .B1 (n_1947),
       .C0 (n_730), .C1 (n_538), .Y (n_2224));
  OAI222X1 g179577(.A0 (n_772), .A1 (n_662), .B0 (n_642), .B1 (n_1947),
       .C0 (n_765), .C1 (n_538), .Y (n_2223));
  AOI22X1 g179578(.A0 (n_1729), .A1 (n_1186), .B0 (\reg_op1[15]_9652 ),
       .B1 (cpu_state[2]), .Y (n_2222));
  AOI22X1 g179579(.A0 (n_1711), .A1 (n_1176), .B0 (\reg_op1[17]_9654 ),
       .B1 (cpu_state[2]), .Y (n_2221));
  AOI22X1 g179580(.A0 (n_1725), .A1 (n_1177), .B0 (\reg_op1[18]_9655 ),
       .B1 (cpu_state[2]), .Y (n_2220));
  AOI22X1 g179581(.A0 (n_1710), .A1 (n_1182), .B0 (\reg_op1[19]_9656 ),
       .B1 (cpu_state[2]), .Y (n_2219));
  AOI22XL g179582(.A0 (cpu_state[5]), .A1 (n_1730), .B0 (cpu_state[3]),
       .B1 (n_6976), .Y (n_2218));
  AOI22X1 g179583(.A0 (cpu_state[5]), .A1 (n_1717), .B0 (n_967), .B1
       (mem_rdata[28]), .Y (n_2217));
  AOI22X1 g179584(.A0 (reg_op1[0]), .A1 (n_1944), .B0 (reg_pc[4]), .B1
       (n_547), .Y (n_2216));
  AOI22X1 g179585(.A0 (\reg_op1[23]_9660 ), .A1 (n_1944), .B0
       (reg_pc[27]), .B1 (n_547), .Y (n_2215));
  AOI22X1 g179586(.A0 (\reg_op1[1]_9638 ), .A1 (n_1944), .B0
       (reg_pc[5]), .B1 (n_547), .Y (n_2214));
  AOI22X1 g179587(.A0 (\reg_op1[2]_9639 ), .A1 (n_1944), .B0
       (reg_pc[6]), .B1 (n_547), .Y (n_2213));
  AOI22X1 g179588(.A0 (\reg_op1[22]_9659 ), .A1 (n_1944), .B0
       (reg_pc[26]), .B1 (n_547), .Y (n_2212));
  AOI22X1 g179589(.A0 (\reg_op1[4]_9641 ), .A1 (n_1944), .B0
       (reg_pc[8]), .B1 (n_547), .Y (n_2211));
  AOI22X1 g179590(.A0 (\reg_op1[5]_9642 ), .A1 (n_1944), .B0
       (reg_pc[9]), .B1 (n_547), .Y (n_2210));
  AOI22X1 g179591(.A0 (\reg_op1[6]_9643 ), .A1 (n_1944), .B0
       (reg_pc[10]), .B1 (n_547), .Y (n_2209));
  AOI22X1 g179592(.A0 (\reg_op1[7]_9644 ), .A1 (n_1944), .B0
       (reg_pc[11]), .B1 (n_547), .Y (n_2208));
  AOI22X1 g179593(.A0 (\reg_op1[8]_9645 ), .A1 (n_1944), .B0
       (reg_pc[12]), .B1 (n_547), .Y (n_2207));
  AOI22X1 g179594(.A0 (\reg_op1[9]_9646 ), .A1 (n_1944), .B0
       (reg_pc[13]), .B1 (n_547), .Y (n_2206));
  AOI22XL g179595(.A0 (\reg_op1[4]_9641 ), .A1 (n_332), .B0 (n_6960),
       .B1 (n_833), .Y (n_2205));
  AOI22X1 g179596(.A0 (\reg_op1[11]_9648 ), .A1 (n_1944), .B0
       (reg_pc[15]), .B1 (n_547), .Y (n_2204));
  AOI22XL g179597(.A0 (\reg_op1[15]_9652 ), .A1 (n_1941), .B0 (n_833),
       .B1 (n_6944), .Y (n_2203));
  AOI22X1 g179598(.A0 (\reg_op1[13]_9650 ), .A1 (n_1944), .B0
       (reg_pc[17]), .B1 (n_547), .Y (n_2202));
  AOI22X1 g179599(.A0 (\reg_op1[22]_9659 ), .A1 (n_550), .B0
       (reg_pc[21]), .B1 (n_547), .Y (n_2201));
  AOI22X1 g179600(.A0 (\reg_op1[20]_9657 ), .A1 (n_1944), .B0
       (reg_pc[24]), .B1 (n_547), .Y (n_2200));
  AOI22XL g179601(.A0 (\reg_op1[24]_9661 ), .A1 (n_1941), .B0 (n_833),
       .B1 (n_6935), .Y (n_2199));
  AOI22X1 g179602(.A0 (n_1805), .A1 (n_673), .B0 (decoded_imm_j[9]),
       .B1 (n_953), .Y (n_2198));
  AOI22X1 g179603(.A0 (\reg_op1[25]_9662 ), .A1 (n_1944), .B0
       (reg_pc[29]), .B1 (n_547), .Y (n_2197));
  AOI22XL g179604(.A0 (\reg_op1[28]_9665 ), .A1 (n_1941), .B0 (n_833),
       .B1 (n_6931), .Y (n_2196));
  AOI22X1 g179605(.A0 (cpu_state[5]), .A1 (n_1721), .B0 (n_967), .B1
       (mem_rdata[26]), .Y (n_2195));
  AOI22X1 g179606(.A0 (cpu_state[5]), .A1 (n_1718), .B0 (n_967), .B1
       (mem_rdata[27]), .Y (n_2194));
  AOI22X1 g179607(.A0 (cpu_state[5]), .A1 (n_1719), .B0 (n_967), .B1
       (mem_rdata[29]), .Y (n_2193));
  AOI22X1 g179608(.A0 (cpu_state[5]), .A1 (n_1723), .B0 (n_967), .B1
       (mem_rdata[30]), .Y (n_2192));
  AOI22XL g179609(.A0 (cpu_state[5]), .A1 (n_1724), .B0 (cpu_state[3]),
       .B1 (n_6985), .Y (n_2191));
  NAND3BXL g179610(.AN (n_6), .B (\reg_op1[8]_9645 ), .C
       (\genblk2.pcpi_div_minus_2470_59_n_492 ), .Y (n_2190));
  NAND4XL g179611(.A (n_985), .B (n_1633), .C (n_305), .D (n_1954), .Y
       (n_2189));
  AOI22X1 g179612(.A0 (\reg_op1[29]_9666 ), .A1 (n_332), .B0
       (\reg_op1[21]_9658 ), .B1 (n_1944), .Y (n_2188));
  OAI22X1 g179613(.A0 (n_717), .A1 (n_677), .B0 (n_577), .B1 (n_1940),
       .Y (n_2187));
  AOI32X1 g179614(.A0 (instr_lb), .A1 (cpu_state[0]), .A2 (n_1949), .B0
       (latched_is_lb), .B1 (n_1948), .Y (n_2186));
  AOI32X1 g179615(.A0 (instr_lh), .A1 (cpu_state[0]), .A2 (n_1949), .B0
       (latched_is_lh), .B1 (n_1948), .Y (n_2185));
  AOI32X1 g179616(.A0 (is_lbu_lhu_lw), .A1 (cpu_state[0]), .A2
       (n_1949), .B0 (latched_is_lu), .B1 (n_1948), .Y (n_2184));
  AOI22X1 g179617(.A0 (\reg_op1[24]_9661 ), .A1 (n_332), .B0
       (\reg_op1[16]_9653 ), .B1 (n_1944), .Y (n_2183));
  NAND4XL g179618(.A (n_756), .B (\genblk2.pcpi_div_minus_2470_59_n_500
       ), .C (\genblk2.pcpi_div_minus_2470_59_n_487 ), .D (n_1418), .Y
       (n_2182));
  AOI22X1 g179619(.A0 (\reg_op1[20]_9657 ), .A1 (n_332), .B0
       (\reg_op1[12]_9649 ), .B1 (n_1944), .Y (n_2181));
  OAI22X1 g179620(.A0 (n_577), .A1 (n_677), .B0 (n_628), .B1 (n_1940),
       .Y (n_2180));
  OAI222X1 g179621(.A0 (n_643), .A1 (n_851), .B0 (n_588), .B1 (n_34),
       .C0 (n_605), .C1 (n_538), .Y (n_2179));
  OAI22X1 g179622(.A0 (n_578), .A1 (n_677), .B0 (n_565), .B1 (n_1940),
       .Y (n_2178));
  AOI22X1 g179623(.A0 (\reg_op1[24]_9661 ), .A1 (n_550), .B0
       (\reg_op1[27]_9664 ), .B1 (n_332), .Y (n_2177));
  INVX1 g179625(.A (n_2174), .Y (n_2175));
  INVX1 g179626(.A (n_2162), .Y (n_2163));
  NOR2X1 g179627(.A (n_1755), .B (n_544), .Y (n_2161));
  NAND2X1 g179629(.A (\reg_op1[6]_9643 ), .B (n_1941), .Y (n_2159));
  NAND2X1 g179630(.A (\reg_op1[24]_9661 ), .B (n_1944), .Y (n_2158));
  OR4X1 g179632(.A (\genblk2.pcpi_div_quotient_msk [10]), .B
       (\genblk2.pcpi_div_quotient_msk [9]), .C
       (\genblk2.pcpi_div_quotient_msk [8]), .D (n_1231), .Y (n_2157));
  NOR4X1 g179633(.A (latched_is_lb), .B (n_931), .C (n_1300), .D
       (n_990), .Y (n_2156));
  OR2X1 g179728(.A (n_1815), .B (n_342), .Y (n_2176));
  NAND2X1 g179730(.A (n_1813), .B (n_673), .Y (n_2174));
  NAND2X1 g179732(.A (n_1811), .B (n_673), .Y (n_2173));
  NAND2X1 g179733(.A (n_1810), .B (n_673), .Y (n_2172));
  NAND2X1 g179734(.A (n_1812), .B (n_673), .Y (n_2171));
  OR2X1 g179735(.A (n_1807), .B (n_342), .Y (n_2170));
  NOR2X1 g179736(.A (n_1803), .B (n_342), .Y (n_2169));
  OR2X1 g179738(.A (n_1958), .B (n_342), .Y (n_2168));
  OR2X1 g179739(.A (n_1802), .B (n_342), .Y (n_2167));
  NOR2X1 g179740(.A (n_850), .B (n_1953), .Y (n_2155));
  NOR2X1 g179742(.A (n_850), .B (n_293), .Y (n_2154));
  NOR2X1 g179743(.A (n_293), .B (n_1953), .Y (n_2166));
  NAND2X1 g179810(.A (cpu_state[2]), .B (n_1955), .Y (n_2165));
  NOR2X1 g179816(.A (n_564), .B (n_1951), .Y (n_2164));
  NOR2X1 g179817(.A (n_636), .B (n_1947), .Y (n_2162));
  INVX1 g179819(.A (n_2146), .Y (n_2145));
  INVX1 g179820(.A (n_2144), .Y (n_2143));
  INVX1 g179831(.A (n_317), .Y (n_2131));
  NAND4XL g179833(.A (n_1153), .B (n_1076), .C (n_1560), .D (n_1100),
       .Y (n_2128));
  OAI21X1 g179834(.A0 (n_1358), .A1 (n_1421), .B0 (n_1541), .Y
       (n_2127));
  OAI21X1 g179835(.A0 (n_622), .A1 (n_1634), .B0 (n_723), .Y (n_2126));
  OAI21X1 g179836(.A0 (n_562), .A1 (n_1630), .B0 (n_1632), .Y (n_2125));
  OAI2BB1X1 g179837(.A0N (n_851), .A1N (n_34), .B0 (mem_rdata_q[31]),
       .Y (n_2124));
  OAI2BB1X1 g179838(.A0N (n_1556), .A1N (n_1637), .B0
       (\reg_op1[31]_9668 ), .Y (n_2123));
  OAI211X1 g179839(.A0 (n_809), .A1 (n_119), .B0 (n_1546), .C0
       (n_1410), .Y (n_2122));
  OAI211X1 g179840(.A0 (n_791), .A1 (n_119), .B0 (n_1548), .C0
       (n_1409), .Y (n_2121));
  OAI221X1 g179841(.A0 (n_278), .A1 (n_1352), .B0 (n_937), .B1 (n_119),
       .C0 (n_1407), .Y (n_2120));
  OAI221X1 g179842(.A0 (n_278), .A1 (n_1359), .B0 (n_897), .B1 (n_119),
       .C0 (n_1415), .Y (n_2119));
  OAI221X1 g179843(.A0 (n_278), .A1 (n_1360), .B0 (n_914), .B1 (n_119),
       .C0 (n_1414), .Y (n_2118));
  OAI211X1 g179844(.A0 (n_803), .A1 (n_119), .B0 (n_1542), .C0
       (n_1413), .Y (n_2117));
  OAI211X1 g179845(.A0 (n_900), .A1 (n_119), .B0 (n_1547), .C0
       (n_1406), .Y (n_2116));
  OAI211X1 g179846(.A0 (n_940), .A1 (n_119), .B0 (n_1545), .C0
       (n_1419), .Y (n_2115));
  OAI221X1 g179847(.A0 (n_278), .A1 (n_1349), .B0 (n_785), .B1 (n_119),
       .C0 (n_1417), .Y (n_2114));
  AOI32X1 g179848(.A0 (\reg_op1[9]_9646 ), .A1 (n_714), .A2 (n_1350),
       .B0 (n_5), .B1 (n_1307), .Y (n_2113));
  AOI22X1 g179850(.A0 (cpu_state[2]), .A1 (n_1629), .B0 (reg_sh[0]),
       .B1 (n_1631), .Y (n_2111));
  AOI22X1 g179851(.A0 (\cpuregs[9] [1]), .A1 (n_1591), .B0
       (\cpuregs[10] [1]), .B1 (n_1601), .Y (n_2110));
  AOI22XL g179852(.A0 (n_434), .A1 (\genblk2.pcpi_div_n_2010 ), .B0
       (\reg_op2[19]_9688 ), .B1 (n_1584), .Y (n_2109));
  AOI22XL g179853(.A0 (n_434), .A1 (\genblk2.pcpi_div_n_2008 ), .B0
       (\reg_op2[21]_9690 ), .B1 (n_1584), .Y (n_2108));
  AOI22XL g179854(.A0 (n_434), .A1 (\genblk2.pcpi_div_n_2007 ), .B0
       (\reg_op2[22]_9691 ), .B1 (n_1584), .Y (n_2107));
  AOI22XL g179855(.A0 (n_434), .A1 (\genblk2.pcpi_div_n_2006 ), .B0
       (\reg_op2[23]_9692 ), .B1 (n_1584), .Y (n_2106));
  AOI22XL g179856(.A0 (n_434), .A1 (\genblk2.pcpi_div_n_1999 ), .B0
       (\reg_op2[30]_9699 ), .B1 (n_1584), .Y (n_2105));
  OAI2BB1X1 g179857(.A0N (n_5692), .A1N (n_1341), .B0 (n_1873), .Y
       (n_2104));
  AOI22X1 g179858(.A0 (reg_next_pc[1]), .A1 (n_1586), .B0 (n_160), .B1
       (n_436), .Y (n_2103));
  AOI22X1 g179859(.A0 (reg_next_pc[2]), .A1 (n_1586), .B0 (n_166), .B1
       (n_436), .Y (n_2102));
  AOI22X1 g179860(.A0 (reg_next_pc[3]), .A1 (n_1586), .B0 (n_168), .B1
       (n_436), .Y (n_2101));
  AOI22X1 g179861(.A0 (reg_next_pc[4]), .A1 (n_1586), .B0 (n_170), .B1
       (n_436), .Y (n_2100));
  AOI22X1 g179862(.A0 (reg_next_pc[5]), .A1 (n_1586), .B0 (n_164), .B1
       (n_436), .Y (n_2099));
  AOI22X1 g179863(.A0 (reg_next_pc[6]), .A1 (n_1586), .B0 (n_174), .B1
       (n_436), .Y (n_2098));
  AOI22X1 g179864(.A0 (reg_next_pc[7]), .A1 (n_1586), .B0 (n_176), .B1
       (n_436), .Y (n_2097));
  AOI22X1 g179865(.A0 (reg_next_pc[8]), .A1 (n_1586), .B0 (n_178), .B1
       (n_436), .Y (n_2096));
  AOI22X1 g179866(.A0 (reg_next_pc[9]), .A1 (n_1586), .B0 (n_180), .B1
       (n_436), .Y (n_2095));
  AOI22X1 g179867(.A0 (reg_next_pc[10]), .A1 (n_1586), .B0 (n_182), .B1
       (n_436), .Y (n_2094));
  AOI22X1 g179868(.A0 (reg_next_pc[11]), .A1 (n_1586), .B0 (n_184), .B1
       (n_436), .Y (n_2093));
  AOI22X1 g179869(.A0 (reg_next_pc[12]), .A1 (n_1586), .B0 (n_186), .B1
       (n_436), .Y (n_2092));
  AOI22X1 g179870(.A0 (reg_next_pc[13]), .A1 (n_1586), .B0 (n_172), .B1
       (n_436), .Y (n_2091));
  AOI22X1 g179871(.A0 (reg_next_pc[14]), .A1 (n_1586), .B0 (n_188), .B1
       (n_436), .Y (n_2090));
  AOI22X1 g179872(.A0 (reg_next_pc[15]), .A1 (n_1586), .B0 (n_190), .B1
       (n_436), .Y (n_2089));
  AOI22X1 g179873(.A0 (reg_next_pc[16]), .A1 (n_1586), .B0 (n_192), .B1
       (n_436), .Y (n_2088));
  AOI22X1 g179874(.A0 (reg_next_pc[17]), .A1 (n_1586), .B0 (n_194), .B1
       (n_436), .Y (n_2087));
  AOI22X1 g179875(.A0 (reg_next_pc[18]), .A1 (n_1586), .B0 (n_196), .B1
       (n_436), .Y (n_2086));
  AOI22X1 g179876(.A0 (reg_next_pc[19]), .A1 (n_1586), .B0 (n_142), .B1
       (n_436), .Y (n_2085));
  AOI22X1 g179877(.A0 (reg_next_pc[20]), .A1 (n_1586), .B0 (n_198), .B1
       (n_436), .Y (n_2084));
  AOI22X1 g179878(.A0 (reg_next_pc[21]), .A1 (n_1586), .B0 (n_144), .B1
       (n_436), .Y (n_2083));
  AOI22X1 g179879(.A0 (reg_next_pc[22]), .A1 (n_1586), .B0 (n_146), .B1
       (n_436), .Y (n_2082));
  AOI22X1 g179880(.A0 (reg_next_pc[23]), .A1 (n_1586), .B0 (n_200), .B1
       (n_436), .Y (n_2081));
  AOI22X1 g179881(.A0 (reg_next_pc[24]), .A1 (n_1586), .B0 (n_202), .B1
       (n_436), .Y (n_2080));
  AOI22X1 g179882(.A0 (reg_next_pc[25]), .A1 (n_1586), .B0 (n_204), .B1
       (n_436), .Y (n_2079));
  AOI22X1 g179883(.A0 (reg_next_pc[26]), .A1 (n_1586), .B0 (n_206), .B1
       (n_436), .Y (n_2078));
  AOI22X1 g179884(.A0 (reg_next_pc[27]), .A1 (n_1586), .B0 (n_208), .B1
       (n_436), .Y (n_2077));
  AOI22X1 g179885(.A0 (reg_next_pc[28]), .A1 (n_1586), .B0 (n_210), .B1
       (n_436), .Y (n_2076));
  AOI22X1 g179886(.A0 (reg_next_pc[29]), .A1 (n_1586), .B0 (n_212), .B1
       (n_436), .Y (n_2075));
  AOI22X1 g179887(.A0 (reg_next_pc[30]), .A1 (n_1586), .B0 (n_214), .B1
       (n_436), .Y (n_2074));
  AOI22X1 g179888(.A0 (reg_next_pc[31]), .A1 (n_1586), .B0 (n_216), .B1
       (n_436), .Y (n_2073));
  AOI22X1 g179889(.A0 (\cpuregs[20] [4]), .A1 (n_1616), .B0
       (\cpuregs[21] [4]), .B1 (n_1614), .Y (n_2072));
  AOI22X1 g179890(.A0 (\cpuregs[28] [4]), .A1 (n_9), .B0
       (\cpuregs[29] [4]), .B1 (n_1599), .Y (n_2071));
  AOI22X1 g179891(.A0 (\cpuregs[24] [0]), .A1 (n_1604), .B0
       (\cpuregs[31] [0]), .B1 (n_1592), .Y (n_2070));
  AOI22X1 g179892(.A0 (\cpuregs[12] [4]), .A1 (n_1610), .B0
       (\cpuregs[11] [4]), .B1 (n_1608), .Y (n_2069));
  AOI22X1 g179893(.A0 (\cpuregs[4] [4]), .A1 (n_1618), .B0
       (\cpuregs[15] [4]), .B1 (n_1593), .Y (n_2068));
  AOI22X1 g179894(.A0 (\cpuregs[12] [2]), .A1 (n_1610), .B0
       (\cpuregs[11] [2]), .B1 (n_1608), .Y (n_2067));
  AOI22X1 g179895(.A0 (\cpuregs[5] [4]), .A1 (n_1611), .B0
       (\cpuregs[6] [4]), .B1 (n_1624), .Y (n_2066));
  AOI22X1 g179896(.A0 (\cpuregs[16] [3]), .A1 (n_1596), .B0
       (\cpuregs[17] [3]), .B1 (n_1625), .Y (n_2065));
  AOI22X1 g179897(.A0 (\cpuregs[4] [3]), .A1 (n_1618), .B0
       (\cpuregs[3] [3]), .B1 (n_1607), .Y (n_2064));
  AOI22X1 g179898(.A0 (\cpuregs[13] [3]), .A1 (n_1606), .B0
       (\cpuregs[14] [3]), .B1 (n_1597), .Y (n_2063));
  AOI22X1 g179899(.A0 (\cpuregs[20] [2]), .A1 (n_1616), .B0
       (\cpuregs[21] [2]), .B1 (n_1614), .Y (n_2062));
  AOI22X1 g179900(.A0 (\cpuregs[24] [2]), .A1 (n_1604), .B0
       (\cpuregs[25] [2]), .B1 (n_1594), .Y (n_2061));
  AOI22X1 g179901(.A0 (\cpuregs[28] [2]), .A1 (n_9), .B0
       (\cpuregs[29] [2]), .B1 (n_1599), .Y (n_2060));
  AOI22X1 g179902(.A0 (\cpuregs[30] [1]), .A1 (n_1622), .B0
       (\cpuregs[31] [1]), .B1 (n_1592), .Y (n_2059));
  AOI22X1 g179903(.A0 (\cpuregs[12] [1]), .A1 (n_1610), .B0
       (\cpuregs[11] [1]), .B1 (n_1608), .Y (n_2058));
  AOI22X1 g179904(.A0 (\cpuregs[8] [1]), .A1 (n_1595), .B0
       (\cpuregs[7] [1]), .B1 (n_1602), .Y (n_2057));
  AOI22X1 g179905(.A0 (\cpuregs[24] [1]), .A1 (n_1604), .B0
       (\cpuregs[25] [1]), .B1 (n_1594), .Y (n_2056));
  AOI22X1 g179906(.A0 (\cpuregs[8] [3]), .A1 (n_1595), .B0
       (\cpuregs[7] [3]), .B1 (n_1602), .Y (n_2055));
  AOI22X1 g179907(.A0 (\cpuregs[9] [0]), .A1 (n_1591), .B0
       (\cpuregs[10] [0]), .B1 (n_1601), .Y (n_2054));
  AOI22X1 g179908(.A0 (\cpuregs[13] [0]), .A1 (n_1606), .B0
       (\cpuregs[14] [0]), .B1 (n_1597), .Y (n_2053));
  AOI22X1 g179909(.A0 (\cpuregs[22] [0]), .A1 (n_1603), .B0
       (\cpuregs[23] [0]), .B1 (n_1627), .Y (n_2052));
  AOI22X1 g179910(.A0 (\cpuregs[20] [1]), .A1 (n_1616), .B0
       (\cpuregs[19] [1]), .B1 (n_1605), .Y (n_2051));
  AOI22X1 g179911(.A0 (\cpuregs[29] [0]), .A1 (n_1599), .B0
       (\cpuregs[30] [0]), .B1 (n_1622), .Y (n_2050));
  AOI22X1 g179913(.A0 (\cpuregs[20] [0]), .A1 (n_1616), .B0
       (\cpuregs[21] [0]), .B1 (n_1614), .Y (n_2048));
  AOI22X1 g179914(.A0 (\cpuregs[18] [0]), .A1 (n_10), .B0
       (\cpuregs[19] [0]), .B1 (n_1605), .Y (n_2047));
  AOI22X1 g179915(.A0 (\cpuregs[16] [0]), .A1 (n_1596), .B0
       (\cpuregs[17] [0]), .B1 (n_1625), .Y (n_2046));
  AOI22X1 g179916(.A0 (\cpuregs[4] [0]), .A1 (n_1618), .B0
       (\cpuregs[3] [0]), .B1 (n_1607), .Y (n_2045));
  AOI22X1 g179917(.A0 (\cpuregs[2] [0]), .A1 (n_1621), .B0
       (\cpuregs[6] [0]), .B1 (n_1624), .Y (n_2044));
  AOI22X1 g179918(.A0 (\cpuregs[8] [0]), .A1 (n_1595), .B0
       (\cpuregs[7] [0]), .B1 (n_1602), .Y (n_2043));
  AOI22X1 g179919(.A0 (\cpuregs[12] [0]), .A1 (n_1610), .B0
       (\cpuregs[11] [0]), .B1 (n_1608), .Y (n_2042));
  AOI22X1 g179920(.A0 (\cpuregs[16] [1]), .A1 (n_1596), .B0
       (\cpuregs[21] [1]), .B1 (n_1614), .Y (n_2041));
  AO22X1 g179921(.A0 (\cpuregs[17] [1]), .A1 (n_1625), .B0
       (\cpuregs[22] [1]), .B1 (n_1603), .Y (n_2040));
  AOI22X1 g179922(.A0 (\cpuregs[26] [1]), .A1 (n_1613), .B0
       (\cpuregs[27] [1]), .B1 (n_1598), .Y (n_2039));
  AOI22X1 g179923(.A0 (\cpuregs[28] [1]), .A1 (n_9), .B0
       (\cpuregs[29] [1]), .B1 (n_1599), .Y (n_2038));
  AOI22X1 g179924(.A0 (\cpuregs[4] [1]), .A1 (n_1618), .B0
       (\cpuregs[3] [1]), .B1 (n_1607), .Y (n_2037));
  AOI22X1 g179925(.A0 (\cpuregs[1] [1]), .A1 (n_1626), .B0
       (\cpuregs[6] [1]), .B1 (n_1624), .Y (n_2036));
  AOI22X1 g179926(.A0 (\cpuregs[13] [1]), .A1 (n_1606), .B0
       (\cpuregs[14] [1]), .B1 (n_1597), .Y (n_2035));
  AOI22X1 g179927(.A0 (\cpuregs[4] [2]), .A1 (n_1618), .B0
       (\cpuregs[3] [2]), .B1 (n_1607), .Y (n_2034));
  AOI22X1 g179928(.A0 (\cpuregs[2] [2]), .A1 (n_1621), .B0
       (\cpuregs[6] [2]), .B1 (n_1624), .Y (n_2033));
  AOI22X1 g179929(.A0 (\cpuregs[13] [2]), .A1 (n_1606), .B0
       (\cpuregs[14] [2]), .B1 (n_1597), .Y (n_2032));
  AOI22X1 g179930(.A0 (\cpuregs[8] [2]), .A1 (n_1595), .B0
       (\cpuregs[7] [2]), .B1 (n_1602), .Y (n_2031));
  AOI22X1 g179931(.A0 (\cpuregs[9] [2]), .A1 (n_1591), .B0
       (\cpuregs[10] [2]), .B1 (n_1601), .Y (n_2030));
  AOI22X1 g179932(.A0 (\cpuregs[26] [2]), .A1 (n_1613), .B0
       (\cpuregs[27] [2]), .B1 (n_1598), .Y (n_2029));
  AO22X1 g179933(.A0 (\cpuregs[18] [2]), .A1 (n_10), .B0
       (\cpuregs[19] [2]), .B1 (n_1605), .Y (n_2028));
  AOI22X1 g179934(.A0 (\cpuregs[16] [2]), .A1 (n_1596), .B0
       (\cpuregs[17] [2]), .B1 (n_1625), .Y (n_2027));
  AOI22X1 g179935(.A0 (\cpuregs[2] [3]), .A1 (n_1621), .B0
       (\cpuregs[6] [3]), .B1 (n_1624), .Y (n_2026));
  AOI22X1 g179936(.A0 (\cpuregs[12] [3]), .A1 (n_1610), .B0
       (\cpuregs[11] [3]), .B1 (n_1608), .Y (n_2025));
  AOI22X1 g179937(.A0 (\cpuregs[9] [3]), .A1 (n_1591), .B0
       (\cpuregs[10] [3]), .B1 (n_1601), .Y (n_2024));
  AOI22X1 g179938(.A0 (\cpuregs[18] [3]), .A1 (n_10), .B0
       (\cpuregs[19] [3]), .B1 (n_1605), .Y (n_2023));
  AOI22X1 g179939(.A0 (\cpuregs[20] [3]), .A1 (n_1616), .B0
       (\cpuregs[21] [3]), .B1 (n_1614), .Y (n_2022));
  AOI22X1 g179940(.A0 (\cpuregs[30] [3]), .A1 (n_1622), .B0
       (\cpuregs[31] [3]), .B1 (n_1592), .Y (n_2021));
  AOI22X1 g179941(.A0 (\cpuregs[26] [3]), .A1 (n_1613), .B0
       (\cpuregs[27] [3]), .B1 (n_1598), .Y (n_2020));
  AO22X1 g179942(.A0 (\cpuregs[24] [3]), .A1 (n_1604), .B0
       (\cpuregs[25] [3]), .B1 (n_1594), .Y (n_2019));
  AOI22X1 g179943(.A0 (\cpuregs[2] [4]), .A1 (n_1621), .B0
       (\cpuregs[3] [4]), .B1 (n_1607), .Y (n_2018));
  AOI22X1 g179944(.A0 (\cpuregs[13] [4]), .A1 (n_1606), .B0
       (\cpuregs[14] [4]), .B1 (n_1597), .Y (n_2017));
  AOI22X1 g179945(.A0 (\cpuregs[8] [4]), .A1 (n_1595), .B0
       (\cpuregs[7] [4]), .B1 (n_1602), .Y (n_2016));
  AOI22X1 g179946(.A0 (\cpuregs[9] [4]), .A1 (n_1591), .B0
       (\cpuregs[10] [4]), .B1 (n_1601), .Y (n_2015));
  AOI22X1 g179947(.A0 (\cpuregs[24] [4]), .A1 (n_1604), .B0
       (\cpuregs[25] [4]), .B1 (n_1594), .Y (n_2014));
  AOI22X1 g179948(.A0 (\cpuregs[26] [4]), .A1 (n_1613), .B0
       (\cpuregs[27] [4]), .B1 (n_1598), .Y (n_2013));
  AOI22X1 g179949(.A0 (\cpuregs[18] [4]), .A1 (n_10), .B0
       (\cpuregs[19] [4]), .B1 (n_1605), .Y (n_2012));
  AO22X1 g179950(.A0 (\cpuregs[16] [4]), .A1 (n_1596), .B0
       (\cpuregs[17] [4]), .B1 (n_1625), .Y (n_2011));
  OAI22X1 g179951(.A0 (n_573), .A1 (n_1637), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_172 ), .B1 (n_1310), .Y
       (n_2010));
  MX2X1 g179952(.A (instr_jalr), .B (n_595), .S0 (n_1357), .Y (n_2009));
  AOI32X1 g179964(.A0 (is_beq_bne_blt_bge_bltu_bgeu), .A1 (n_538), .A2
       (n_1321), .B0 (instr_bne), .B1 (n_537), .Y (n_1997));
  OAI2BB1X1 g179965(.A0N (instr_lh), .A1N (n_537), .B0 (n_1929), .Y
       (n_1996));
  OAI2BB1X1 g179966(.A0N (instr_sh), .A1N (n_537), .B0 (n_1928), .Y
       (n_1995));
  AOI32X1 g179967(.A0 (is_alu_reg_imm), .A1 (n_538), .A2 (n_1323), .B0
       (instr_addi), .B1 (n_537), .Y (n_1994));
  AOI32X1 g179968(.A0 (is_beq_bne_blt_bge_bltu_bgeu), .A1 (n_538), .A2
       (n_1323), .B0 (instr_beq), .B1 (n_537), .Y (n_1993));
  OAI2BB1X1 g179969(.A0N (instr_lb), .A1N (n_537), .B0 (n_1927), .Y
       (n_1992));
  OAI2BB1X1 g179970(.A0N (instr_sb), .A1N (n_537), .B0 (n_1925), .Y
       (n_1991));
  OAI2BB1X1 g179971(.A0N (instr_lhu), .A1N (n_537), .B0 (n_1926), .Y
       (n_1990));
  AOI32X1 g179972(.A0 (is_beq_bne_blt_bge_bltu_bgeu), .A1 (n_538), .A2
       (n_1325), .B0 (instr_bge), .B1 (n_537), .Y (n_1989));
  AOI32X1 g179973(.A0 (is_alu_reg_imm), .A1 (n_538), .A2 (n_1338), .B0
       (instr_andi), .B1 (n_537), .Y (n_1988));
  AOI32X1 g179974(.A0 (is_beq_bne_blt_bge_bltu_bgeu), .A1 (n_538), .A2
       (n_1338), .B0 (instr_bgeu), .B1 (n_537), .Y (n_1987));
  AOI32X1 g179975(.A0 (is_beq_bne_blt_bge_bltu_bgeu), .A1 (n_538), .A2
       (n_1337), .B0 (instr_blt), .B1 (n_537), .Y (n_1986));
  AOI32X1 g179976(.A0 (is_beq_bne_blt_bge_bltu_bgeu), .A1 (n_538), .A2
       (n_1344), .B0 (instr_bltu), .B1 (n_537), .Y (n_1985));
  OAI2BB1X1 g179977(.A0N (instr_lbu), .A1N (n_537), .B0 (n_1923), .Y
       (n_1984));
  OAI2BB1X1 g179978(.A0N (instr_lw), .A1N (n_537), .B0 (n_1924), .Y
       (n_1983));
  AOI32X1 g179979(.A0 (is_alu_reg_imm), .A1 (n_538), .A2 (n_1344), .B0
       (instr_ori), .B1 (n_537), .Y (n_1982));
  AOI32X1 g179980(.A0 (is_alu_reg_imm), .A1 (n_538), .A2 (n_1326), .B0
       (instr_slti), .B1 (n_537), .Y (n_1981));
  OAI2BB1X1 g179981(.A0N (instr_sw), .A1N (n_537), .B0 (n_1922), .Y
       (n_1980));
  AOI32X1 g179982(.A0 (is_alu_reg_imm), .A1 (n_538), .A2 (n_1337), .B0
       (instr_xori), .B1 (n_537), .Y (n_1979));
  OAI32X1 g179984(.A0 (latched_rd[0]), .A1 (latched_rd[3]), .A2
       (n_1331), .B0 (latched_branch), .B1 (n_442), .Y (n_1977));
  NOR4X1 g179985(.A (mem_rdata_q[4]), .B (mem_rdata_q[5]), .C
       (mem_rdata_q[0]), .D (n_1215), .Y (n_1976));
  AOI32X1 g179987(.A0 (\reg_op2[1]_9670 ), .A1 (\reg_op1[1]_9638 ), .A2
       (n_283), .B0 (is_lui_auipc_jal_jalr_addi_add_sub), .B1 (n_6626),
       .Y (n_1974));
  NOR3X1 g180003(.A (mem_rdata_q[31]), .B (n_579), .C (n_1639), .Y
       (n_2153));
  AOI31X1 g180004(.A0 (n_562), .A1 (mem_rdata[1]), .A2 (mem_rdata[0]),
       .B0 (n_1957), .Y (n_2152));
  NOR2X1 g180005(.A (n_1525), .B (n_1955), .Y (n_2151));
  NOR3X1 g180006(.A (n_6554), .B (n_60), .C (n_1950), .Y (n_2150));
  NAND3X1 g180007(.A (n_288), .B (n_356), .C (n_1633), .Y (n_305));
  NOR3X1 g180008(.A (mem_rdata_q[31]), .B (mem_rdata_q[30]), .C
       (n_1639), .Y (n_323));
  OAI211X1 g180009(.A0 (n_277), .A1 (n_1213), .B0 (n_821), .C0
       (n_1029), .Y (n_326));
  OAI211X1 g180010(.A0 (n_277), .A1 (n_1212), .B0 (n_935), .C0
       (n_1035), .Y (n_2146));
  OAI211X1 g180011(.A0 (n_277), .A1 (n_1210), .B0 (n_786), .C0
       (n_1034), .Y (n_2144));
  OAI221X1 g180012(.A0 (n_268), .A1 (n_1204), .B0 (n_277), .B1
       (n_1201), .C0 (n_892), .Y (n_439));
  OAI211X1 g180013(.A0 (n_277), .A1 (n_1200), .B0 (n_810), .C0
       (n_1081), .Y (n_327));
  OAI211X1 g180014(.A0 (n_277), .A1 (n_1211), .B0 (n_930), .C0
       (n_1036), .Y (n_2140));
  OAI221X1 g180015(.A0 (n_268), .A1 (n_1197), .B0 (n_277), .B1
       (n_1208), .C0 (n_915), .Y (n_438));
  NAND2X1 g180016(.A (n_1033), .B (n_1799), .Y (n_503));
  OAI211X1 g180017(.A0 (n_277), .A1 (n_1206), .B0 (n_788), .C0
       (n_1031), .Y (n_2137));
  OAI221X1 g180018(.A0 (n_277), .A1 (n_1214), .B0 (n_268), .B1
       (n_1362), .C0 (n_921), .Y (n_437));
  NAND2X1 g180019(.A (n_1032), .B (n_1798), .Y (n_440));
  OAI211X1 g180020(.A0 (n_277), .A1 (n_1209), .B0 (n_823), .C0
       (n_1037), .Y (n_504));
  OAI211X1 g180021(.A0 (n_277), .A1 (n_1202), .B0 (n_824), .C0
       (n_1030), .Y (n_334));
  NAND2X1 g180022(.A (n_1028), .B (n_1937), .Y (n_317));
  AO22X2 g180023(.A0 (n_555), .A1 (n_1536), .B0 (reg_out[0]), .B1
       (n_11742), .Y (n_358));
  INVX1 g180024(.A (n_1949), .Y (n_1948));
  INVX1 g180025(.A (n_1947), .Y (n_1946));
  INVX1 g180027(.A (n_1944), .Y (n_1943));
  INVX1 g180029(.A (n_1941), .Y (n_1940));
  AOI222X1 g180030(.A0 (n_971), .A1 (mem_rdata[12]), .B0 (n_970), .B1
       (mem_rdata[20]), .C0 (\reg_op1[4]_9641 ), .C1 (cpu_state[2]), .Y
       (n_1939));
  AOI222X1 g180031(.A0 (n_971), .A1 (mem_rdata[10]), .B0 (n_970), .B1
       (mem_rdata[18]), .C0 (\reg_op1[2]_9639 ), .C1 (cpu_state[2]), .Y
       (n_1938));
  AOI22X1 g180032(.A0 (n_567), .A1 (n_1207), .B0
       (mem_16bit_buffer[12]), .B1 (n_360), .Y (n_1937));
  AOI21X1 g180034(.A0 (n_2), .A1 (n_50), .B0 (cpu_state[5]), .Y
       (n_1935));
  OAI2BB1X1 g180035(.A0N (n_2), .A1N (n_114), .B0 (n_548), .Y (n_1934));
  OAI2BB1X1 g180036(.A0N (n_2), .A1N (n_64), .B0 (n_548), .Y (n_1933));
  OAI2BB1X1 g180037(.A0N (n_2), .A1N (n_62), .B0 (n_548), .Y (n_1932));
  OAI2BB1X1 g180038(.A0N (n_2), .A1N (n_66), .B0 (n_548), .Y (n_1931));
  OAI2BB1X1 g180039(.A0N (n_2), .A1N (n_68), .B0 (n_548), .Y (n_1930));
  NAND3X1 g180040(.A (is_lb_lh_lw_lbu_lhu), .B (n_538), .C (n_1321), .Y
       (n_1929));
  NAND3X1 g180041(.A (is_sb_sh_sw), .B (n_538), .C (n_1321), .Y
       (n_1928));
  NAND3X1 g180042(.A (is_lb_lh_lw_lbu_lhu), .B (n_538), .C (n_1323), .Y
       (n_1927));
  NAND3X1 g180043(.A (is_lb_lh_lw_lbu_lhu), .B (n_538), .C (n_1325), .Y
       (n_1926));
  NAND3X1 g180044(.A (is_sb_sh_sw), .B (n_538), .C (n_1323), .Y
       (n_1925));
  NAND3X1 g180045(.A (is_lb_lh_lw_lbu_lhu), .B (n_538), .C (n_1326), .Y
       (n_1924));
  NAND3X1 g180046(.A (is_lb_lh_lw_lbu_lhu), .B (n_538), .C (n_1337), .Y
       (n_1923));
  NAND3X1 g180047(.A (is_sb_sh_sw), .B (n_538), .C (n_1326), .Y
       (n_1922));
  AOI21XL g180048(.A0 (n_6543), .A1 (n_1248), .B0 (n_986), .Y (n_1921));
  OAI2BB1X1 g180049(.A0N (n_1302), .A1N (n_258), .B0 (n_307), .Y
       (n_1920));
  OAI2BB1X1 g180050(.A0N (n_1301), .A1N (n_258), .B0 (n_307), .Y
       (n_1919));
  OAI21XL g180051(.A0 (mem_ready), .A1 (n_545), .B0 (n_1630), .Y
       (n_1918));
  NOR2X1 g180052(.A (n_1420), .B (n_544), .Y (n_1917));
  OR2X1 g180053(.A (n_278), .B (n_1194), .Y (n_1916));
  NAND2X1 g180054(.A (n_279), .B (n_1198), .Y (n_1915));
  NOR2X1 g180055(.A (n_565), .B (n_878), .Y (n_1914));
  NOR2X1 g180056(.A (n_544), .B (n_1384), .Y (n_1913));
  NOR2X1 g180057(.A (n_544), .B (n_1405), .Y (n_1912));
  NOR2X1 g180058(.A (n_544), .B (n_1377), .Y (n_1911));
  NOR2X1 g180059(.A (n_544), .B (n_1386), .Y (n_1910));
  NOR2X1 g180060(.A (n_544), .B (n_1452), .Y (n_1909));
  NOR2X1 g180061(.A (n_544), .B (n_1432), .Y (n_1908));
  NOR2X1 g180062(.A (n_544), .B (n_1424), .Y (n_1907));
  NOR2X1 g180063(.A (n_544), .B (n_1474), .Y (n_1906));
  NOR2X1 g180064(.A (n_544), .B (n_1473), .Y (n_1905));
  NOR2X1 g180065(.A (n_544), .B (n_1430), .Y (n_1904));
  NAND2BX1 g180066(.AN (n_1629), .B (reg_sh[1]), .Y (n_1903));
  NOR2X1 g180067(.A (n_1440), .B (n_544), .Y (n_1902));
  NAND2XL g180068(.A (\genblk2.pcpi_div_n_2028 ), .B (n_434), .Y
       (n_1901));
  NAND2XL g180069(.A (\genblk2.pcpi_div_n_2027 ), .B (n_434), .Y
       (n_1900));
  NAND2XL g180070(.A (\genblk2.pcpi_div_n_2026 ), .B (n_434), .Y
       (n_1899));
  NAND2XL g180071(.A (\genblk2.pcpi_div_n_2025 ), .B (n_434), .Y
       (n_1898));
  NAND2XL g180072(.A (\genblk2.pcpi_div_n_2024 ), .B (n_434), .Y
       (n_1897));
  NAND2XL g180073(.A (\genblk2.pcpi_div_n_2023 ), .B (n_434), .Y
       (n_1896));
  NAND2XL g180074(.A (\genblk2.pcpi_div_n_2022 ), .B (n_434), .Y
       (n_1895));
  NAND2XL g180075(.A (\genblk2.pcpi_div_n_2021 ), .B (n_434), .Y
       (n_1894));
  NAND2XL g180076(.A (\genblk2.pcpi_div_n_2020 ), .B (n_434), .Y
       (n_1893));
  NAND2XL g180077(.A (\genblk2.pcpi_div_n_2019 ), .B (n_434), .Y
       (n_1892));
  NAND2XL g180078(.A (n_434), .B (\genblk2.pcpi_div_n_2018 ), .Y
       (n_1891));
  NAND2XL g180079(.A (n_434), .B (\genblk2.pcpi_div_n_2017 ), .Y
       (n_1890));
  NAND2XL g180080(.A (n_434), .B (\genblk2.pcpi_div_n_2016 ), .Y
       (n_1889));
  NAND2XL g180081(.A (n_434), .B (\genblk2.pcpi_div_n_2015 ), .Y
       (n_1888));
  NAND2XL g180082(.A (n_434), .B (\genblk2.pcpi_div_n_2014 ), .Y
       (n_1887));
  NAND2XL g180083(.A (n_434), .B (\genblk2.pcpi_div_n_2013 ), .Y
       (n_1886));
  NOR2X1 g180084(.A (n_544), .B (n_1375), .Y (n_1885));
  NAND2XL g180085(.A (n_434), .B (\genblk2.pcpi_div_n_2012 ), .Y
       (n_1884));
  NAND2XL g180086(.A (n_434), .B (\genblk2.pcpi_div_n_2011 ), .Y
       (n_1883));
  NAND2XL g180087(.A (n_434), .B (\genblk2.pcpi_div_n_2009 ), .Y
       (n_1882));
  NAND2XL g180088(.A (n_434), .B (\genblk2.pcpi_div_n_2005 ), .Y
       (n_1881));
  NAND2XL g180089(.A (n_434), .B (\genblk2.pcpi_div_n_2004 ), .Y
       (n_1880));
  NAND2XL g180090(.A (n_434), .B (\genblk2.pcpi_div_n_2003 ), .Y
       (n_1879));
  NAND2XL g180091(.A (n_434), .B (\genblk2.pcpi_div_n_2002 ), .Y
       (n_1878));
  NAND2XL g180092(.A (n_434), .B (\genblk2.pcpi_div_n_2001 ), .Y
       (n_1877));
  NAND2XL g180093(.A (n_434), .B (\genblk2.pcpi_div_n_2000 ), .Y
       (n_1876));
  NOR2X1 g180094(.A (n_544), .B (n_1372), .Y (n_1875));
  NAND2BX1 g180095(.AN (n_1632), .B (n_48), .Y (n_1874));
  NAND2BX1 g180096(.AN (n_1628), .B (n_313), .Y (n_1873));
  NOR2X1 g180097(.A (n_544), .B (n_1468), .Y (n_1872));
  NAND2BX1 g180098(.AN (n_1628), .B (n_48), .Y (n_1871));
  NOR2X1 g180099(.A (n_544), .B (n_1478), .Y (n_1870));
  NAND2X1 g180100(.A (\cpuregs[1] [4]), .B (n_1626), .Y (n_1869));
  NOR2X1 g180101(.A (n_1466), .B (n_544), .Y (n_1868));
  NAND2X1 g180103(.A (\cpuregs[1] [3]), .B (n_1626), .Y (n_1866));
  NOR2X1 g180104(.A (n_544), .B (n_1470), .Y (n_1865));
  NOR2X1 g180105(.A (n_1444), .B (n_544), .Y (n_1864));
  NAND2X1 g180106(.A (\cpuregs[1] [2]), .B (n_1626), .Y (n_1863));
  OAI2BB1X1 g180107(.A0N (n_545), .A1N (n_804), .B0 (n_1630), .Y
       (n_1862));
  NOR2X1 g180108(.A (n_544), .B (n_1379), .Y (n_1861));
  NOR2X1 g180109(.A (n_544), .B (n_1388), .Y (n_1860));
  NOR2X1 g180110(.A (n_544), .B (n_1404), .Y (n_1859));
  NOR2X1 g180111(.A (n_544), .B (n_1380), .Y (n_1858));
  NOR2X1 g180112(.A (n_544), .B (n_1383), .Y (n_1857));
  NOR2X1 g180113(.A (n_544), .B (n_1472), .Y (n_1856));
  NOR2X1 g180114(.A (n_544), .B (n_1453), .Y (n_1855));
  NOR2X1 g180115(.A (n_544), .B (n_1441), .Y (n_1854));
  NOR2X1 g180116(.A (n_544), .B (n_1403), .Y (n_1853));
  NOR2X1 g180117(.A (n_544), .B (n_1457), .Y (n_1852));
  NOR2X1 g180118(.A (n_544), .B (n_1402), .Y (n_1851));
  NOR2X1 g180119(.A (n_544), .B (n_1401), .Y (n_1850));
  NOR2X1 g180120(.A (n_544), .B (n_1400), .Y (n_1849));
  NOR2X1 g180121(.A (n_544), .B (n_1399), .Y (n_1848));
  NOR2X1 g180122(.A (n_544), .B (n_1398), .Y (n_1847));
  NOR2X1 g180123(.A (n_544), .B (n_1397), .Y (n_1846));
  NOR2X1 g180124(.A (n_544), .B (n_1449), .Y (n_1845));
  NOR2X1 g180125(.A (n_544), .B (n_1395), .Y (n_1844));
  NOR2X1 g180126(.A (n_544), .B (n_1396), .Y (n_1843));
  NOR2X1 g180127(.A (n_544), .B (n_1382), .Y (n_1842));
  NOR2X1 g180128(.A (n_544), .B (n_1394), .Y (n_1841));
  NOR2X1 g180129(.A (n_544), .B (n_1393), .Y (n_1840));
  NOR2X1 g180130(.A (n_544), .B (n_1412), .Y (n_1839));
  NOR2X1 g180131(.A (n_544), .B (n_1392), .Y (n_1838));
  NOR2X1 g180132(.A (n_544), .B (n_1391), .Y (n_1837));
  NOR2X1 g180133(.A (n_544), .B (n_1390), .Y (n_1836));
  NOR2X1 g180134(.A (n_544), .B (n_1389), .Y (n_1835));
  NOR2X1 g180135(.A (n_544), .B (n_1387), .Y (n_1834));
  NOR2X1 g180136(.A (n_544), .B (n_1385), .Y (n_1833));
  NOR2X1 g180137(.A (n_544), .B (n_1469), .Y (n_1832));
  NOR2X1 g180138(.A (n_544), .B (n_1374), .Y (n_1831));
  NOR2X1 g180139(.A (n_544), .B (n_1451), .Y (n_1830));
  NOR2X1 g180140(.A (n_544), .B (n_1479), .Y (n_1829));
  NOR2X1 g180141(.A (n_544), .B (n_1461), .Y (n_1828));
  NOR2X1 g180142(.A (n_544), .B (n_1436), .Y (n_1827));
  NOR2X1 g180143(.A (n_1435), .B (n_544), .Y (n_1826));
  NOR2X1 g180144(.A (n_544), .B (n_1480), .Y (n_1825));
  NOR2X1 g180145(.A (n_544), .B (n_1378), .Y (n_1824));
  NOR2X1 g180146(.A (n_544), .B (n_1477), .Y (n_1823));
  NOR2X1 g180147(.A (n_544), .B (n_1475), .Y (n_1822));
  NOR2X1 g180148(.A (n_544), .B (n_1381), .Y (n_1821));
  NOR2X1 g180149(.A (n_544), .B (n_1434), .Y (n_1820));
  NOR2X1 g180150(.A (n_1437), .B (n_544), .Y (n_1819));
  NOR2X1 g180151(.A (n_544), .B (n_1373), .Y (n_1818));
  NOR2X1 g180152(.A (n_544), .B (n_1376), .Y (n_1817));
  AOI222X1 g180154(.A0 (mem_rdata[1]), .A1 (n_839), .B0
       (mem_rdata_q[1]), .B1 (n_505), .C0 (n_562), .C1 (n_6865), .Y
       (n_1958));
  NAND3BXL g180155(.AN (n_1193), .B (n_545), .C (n_150), .Y (n_1957));
  AOI31X1 g180158(.A0 (n_905), .A1 (n_545), .A2 (n_446), .B0 (n_544),
       .Y (n_1956));
  NOR2BX1 g180160(.AN (n_1629), .B (reg_sh[1]), .Y (n_1955));
  NOR2BX1 g180161(.AN (n_288), .B (n_1638), .Y (n_1954));
  NOR2X1 g180164(.A (n_544), .B (n_1636), .Y (n_1953));
  NOR4X1 g180179(.A (mem_do_wdata), .B (n_761), .C (n_544), .D (n_881),
       .Y (n_293));
  NAND2BX1 g180190(.AN (n_1523), .B (latched_is_lb), .Y (n_1951));
  OA21X1 g180198(.A0 (n_158), .A1 (n_664), .B0 (n_472), .Y (n_1950));
  NAND2X1 g180199(.A (n_615), .B (n_1636), .Y (n_1949));
  AND2X1 g180200(.A (n_1327), .B (n_34), .Y (n_1947));
  AND2X2 g180201(.A (n_1363), .B (n_1631), .Y (n_332));
  AND2X1 g180202(.A (n_993), .B (n_1631), .Y (n_1944));
  AND3X1 g180203(.A (cpu_state[2]), .B (n_1322), .C (n_1363), .Y
       (n_550));
  AND2X1 g180204(.A (cpu_state[2]), .B (n_1529), .Y (n_1941));
  NAND4XL g180205(.A (n_1117), .B (n_1120), .C (n_1113), .D (n_1118),
       .Y (n_1801));
  AOI222X1 g180206(.A0 (n_971), .A1 (mem_rdata[11]), .B0 (n_970), .B1
       (mem_rdata[19]), .C0 (\reg_op1[3]_9640 ), .C1 (cpu_state[2]), .Y
       (n_1800));
  AOI22X1 g180207(.A0 (n_567), .A1 (n_1203), .B0
       (mem_16bit_buffer[10]), .B1 (n_360), .Y (n_1799));
  AOI22X1 g180208(.A0 (n_567), .A1 (n_1205), .B0
       (mem_16bit_buffer[11]), .B1 (n_360), .Y (n_1798));
  AOI222X1 g180209(.A0 (n_971), .A1 (mem_rdata[13]), .B0 (n_970), .B1
       (mem_rdata[21]), .C0 (\reg_op1[5]_9642 ), .C1 (cpu_state[2]), .Y
       (n_1797));
  OR4X1 g180210(.A (n_622), .B (n_616), .C (n_853), .D (n_537), .Y
       (n_1796));
  AOI22X1 g180211(.A0 (n_1318), .A1 (mem_rdata[21]), .B0
       (cpu_state[3]), .B1 (n_94), .Y (n_1795));
  AOI22X1 g180212(.A0 (n_1318), .A1 (mem_rdata[28]), .B0
       (cpu_state[3]), .B1 (n_106), .Y (n_1794));
  AOI22X1 g180213(.A0 (n_1318), .A1 (mem_rdata[26]), .B0
       (cpu_state[3]), .B1 (n_104), .Y (n_1793));
  AOI22X1 g180214(.A0 (n_1318), .A1 (mem_rdata[27]), .B0
       (cpu_state[3]), .B1 (n_108), .Y (n_1792));
  AOI22X1 g180215(.A0 (n_1318), .A1 (mem_rdata[25]), .B0
       (cpu_state[3]), .B1 (n_102), .Y (n_1791));
  AOI22X1 g180216(.A0 (n_1318), .A1 (mem_rdata[30]), .B0
       (cpu_state[3]), .B1 (n_112), .Y (n_1790));
  AOI22X1 g180217(.A0 (n_1318), .A1 (mem_rdata[24]), .B0
       (cpu_state[3]), .B1 (n_100), .Y (n_1789));
  AOI22X1 g180218(.A0 (n_1318), .A1 (mem_rdata[18]), .B0
       (cpu_state[3]), .B1 (n_90), .Y (n_1788));
  AOI22X1 g180219(.A0 (n_1318), .A1 (mem_rdata[16]), .B0
       (\reg_op1[16]_9653 ), .B1 (cpu_state[2]), .Y (n_1787));
  AOI22X1 g180220(.A0 (n_1318), .A1 (mem_rdata[17]), .B0
       (cpu_state[3]), .B1 (n_86), .Y (n_1786));
  AOI22X1 g180221(.A0 (n_1318), .A1 (mem_rdata[23]), .B0
       (cpu_state[3]), .B1 (n_98), .Y (n_1785));
  AOI22X1 g180222(.A0 (n_1318), .A1 (mem_rdata[20]), .B0
       (cpu_state[3]), .B1 (n_88), .Y (n_1784));
  AOI22X1 g180223(.A0 (n_1324), .A1 (mem_rdata[30]), .B0 (n_1320), .B1
       (mem_rdata[14]), .Y (n_1783));
  AO22X1 g180224(.A0 (decoded_imm[31]), .A1 (n_421), .B0
       (\reg_op2[31]_9700 ), .B1 (n_832), .Y (n_1782));
  AOI22X1 g180225(.A0 (n_1318), .A1 (mem_rdata[22]), .B0
       (cpu_state[3]), .B1 (n_96), .Y (n_1781));
  AOI22X1 g180226(.A0 (n_1324), .A1 (mem_rdata[29]), .B0 (n_1320), .B1
       (mem_rdata[13]), .Y (n_1780));
  AOI22X1 g180227(.A0 (n_1324), .A1 (mem_rdata[28]), .B0 (n_1320), .B1
       (mem_rdata[12]), .Y (n_1779));
  AO22X1 g180228(.A0 (decoded_imm[15]), .A1 (n_421), .B0
       (\reg_op2[15]_9684 ), .B1 (n_832), .Y (n_1778));
  AOI22X1 g180229(.A0 (n_1324), .A1 (mem_rdata[24]), .B0 (n_1320), .B1
       (mem_rdata[8]), .Y (n_1777));
  AO22X1 g180230(.A0 (decoded_imm[30]), .A1 (n_421), .B0
       (\reg_op2[30]_9699 ), .B1 (n_832), .Y (n_1776));
  AO22X1 g180231(.A0 (decoded_imm[14]), .A1 (n_421), .B0
       (\reg_op2[14]_9683 ), .B1 (n_832), .Y (n_1775));
  AOI22X1 g180232(.A0 (n_976), .A1 (n_1199), .B0 (cpu_state[3]), .B1
       (n_82), .Y (n_1774));
  AO22X1 g180233(.A0 (decoded_imm[8]), .A1 (n_421), .B0
       (\reg_op2[8]_9677 ), .B1 (n_832), .Y (n_1773));
  AOI22X1 g180234(.A0 (n_1324), .A1 (mem_rdata[27]), .B0 (n_1320), .B1
       (mem_rdata[11]), .Y (n_1772));
  AOI22X1 g180235(.A0 (n_1324), .A1 (mem_rdata[26]), .B0 (n_1320), .B1
       (mem_rdata[10]), .Y (n_1771));
  AOI22X1 g180236(.A0 (n_1324), .A1 (mem_rdata[25]), .B0 (n_1320), .B1
       (mem_rdata[9]), .Y (n_1770));
  AO22X1 g180237(.A0 (decoded_imm[12]), .A1 (n_421), .B0
       (\reg_op2[12]_9681 ), .B1 (n_832), .Y (n_1769));
  AOI22X1 g180238(.A0 (n_1318), .A1 (mem_rdata[29]), .B0
       (cpu_state[3]), .B1 (n_110), .Y (n_1768));
  AO22X1 g180239(.A0 (decoded_imm[9]), .A1 (n_421), .B0
       (\reg_op2[9]_9678 ), .B1 (n_832), .Y (n_1767));
  AO22X1 g180240(.A0 (decoded_imm[11]), .A1 (n_421), .B0
       (\reg_op2[11]_9680 ), .B1 (n_832), .Y (n_1766));
  AO22X1 g180241(.A0 (decoded_imm[13]), .A1 (n_421), .B0
       (\reg_op2[13]_9682 ), .B1 (n_832), .Y (n_1765));
  AO22X1 g180242(.A0 (decoded_imm[16]), .A1 (n_421), .B0
       (\reg_op2[16]_9685 ), .B1 (n_832), .Y (n_1764));
  AO22X1 g180243(.A0 (decoded_imm[18]), .A1 (n_421), .B0
       (\reg_op2[18]_9687 ), .B1 (n_832), .Y (n_1763));
  AO22X1 g180244(.A0 (decoded_imm[19]), .A1 (n_421), .B0
       (\reg_op2[19]_9688 ), .B1 (n_832), .Y (n_1762));
  AO22X1 g180245(.A0 (decoded_imm[20]), .A1 (n_421), .B0
       (\reg_op2[20]_9689 ), .B1 (n_832), .Y (n_1761));
  AO22X1 g180246(.A0 (decoded_imm[21]), .A1 (n_421), .B0
       (\reg_op2[21]_9690 ), .B1 (n_832), .Y (n_1760));
  AO22X1 g180247(.A0 (decoded_imm[22]), .A1 (n_421), .B0
       (\reg_op2[22]_9691 ), .B1 (n_832), .Y (n_1759));
  AO22X1 g180248(.A0 (decoded_imm[25]), .A1 (n_421), .B0
       (\reg_op2[25]_9694 ), .B1 (n_832), .Y (n_1758));
  AO22X1 g180249(.A0 (decoded_imm[27]), .A1 (n_421), .B0
       (\reg_op2[27]_9696 ), .B1 (n_832), .Y (n_1757));
  AOI22X1 g180250(.A0 (n_1318), .A1 (mem_rdata[19]), .B0
       (cpu_state[3]), .B1 (n_92), .Y (n_1756));
  MXI2XL g180251(.A (cpu_state[3]), .B (latched_stalu), .S0 (n_1216),
       .Y (n_1755));
  OAI32X1 g180260(.A0 (n_736), .A1 (n_615), .A2 (n_675), .B0 (n_592),
       .B1 (n_1319), .Y (n_1746));
  OAI32X1 g180261(.A0 (n_777), .A1 (n_615), .A2 (n_675), .B0 (n_580),
       .B1 (n_1319), .Y (n_1745));
  OAI2BB1X1 g180262(.A0N (latched_rd[4]), .A1N (n_675), .B0 (n_1554),
       .Y (n_1744));
  OAI2BB1X1 g180263(.A0N (latched_rd[0]), .A1N (n_675), .B0 (n_1552),
       .Y (n_1743));
  OAI32X1 g180264(.A0 (n_740), .A1 (n_615), .A2 (n_675), .B0 (n_638),
       .B1 (n_1319), .Y (n_1742));
  NAND4XL g180267(.A (n_1115), .B (n_1055), .C (n_1051), .D (n_1162),
       .Y (n_1739));
  NAND4XL g180268(.A (n_1149), .B (n_1148), .C (n_1122), .D (n_1161),
       .Y (n_1738));
  NAND4XL g180269(.A (n_1151), .B (n_1156), .C (n_1152), .D (n_1042),
       .Y (n_1737));
  NAND4XL g180270(.A (n_1157), .B (n_1110), .C (n_1059), .D (n_1054),
       .Y (n_1736));
  NAND4XL g180271(.A (n_1077), .B (n_1154), .C (n_1050), .D (n_1038),
       .Y (n_1735));
  NAND4XL g180272(.A (n_1082), .B (n_1114), .C (n_1070), .D (n_1061),
       .Y (n_1734));
  NAND4XL g180273(.A (n_1140), .B (n_1052), .C (n_1144), .D (n_1142),
       .Y (n_1733));
  NAND4XL g180274(.A (n_1066), .B (n_1063), .C (n_1155), .D (n_1049),
       .Y (n_1732));
  NAND4XL g180275(.A (n_1129), .B (n_1068), .C (n_1048), .D (n_1159),
       .Y (n_1731));
  NAND4XL g180276(.A (n_1143), .B (n_1145), .C (n_1091), .D (n_1062),
       .Y (n_1730));
  NAND4XL g180277(.A (n_1098), .B (n_1138), .C (n_1056), .D (n_1106),
       .Y (n_1729));
  NAND4XL g180278(.A (n_1107), .B (n_1141), .C (n_1133), .D (n_1136),
       .Y (n_1728));
  NAND4XL g180279(.A (n_1078), .B (n_1045), .C (n_1044), .D (n_1073),
       .Y (n_1727));
  NAND4XL g180280(.A (n_1134), .B (n_1060), .C (n_1132), .D (n_1160),
       .Y (n_1726));
  NAND4XL g180281(.A (n_1041), .B (n_1116), .C (n_1109), .D (n_1119),
       .Y (n_1725));
  NAND4XL g180282(.A (n_1065), .B (n_1096), .C (n_1095), .D (n_1057),
       .Y (n_1724));
  NAND4XL g180283(.A (n_1089), .B (n_1092), .C (n_1139), .D (n_1093),
       .Y (n_1723));
  NAND4XL g180284(.A (n_1123), .B (n_1121), .C (n_1103), .D (n_1104),
       .Y (n_1722));
  NAND4XL g180285(.A (n_1080), .B (n_1075), .C (n_1192), .D (n_1158),
       .Y (n_1721));
  NAND4XL g180286(.A (n_1112), .B (n_1099), .C (n_1067), .D (n_1127),
       .Y (n_1720));
  NAND4XL g180287(.A (n_1074), .B (n_1079), .C (n_1088), .D (n_1090),
       .Y (n_1719));
  NAND4XL g180288(.A (n_1083), .B (n_1072), .C (n_1102), .D (n_1084),
       .Y (n_1718));
  NAND4XL g180289(.A (n_1087), .B (n_1137), .C (n_1058), .D (n_1135),
       .Y (n_1717));
  NAND4XL g180290(.A (n_1085), .B (n_1150), .C (n_1097), .D (n_1111),
       .Y (n_1716));
  NAND4XL g180291(.A (n_1086), .B (n_1069), .C (n_1043), .D (n_1047),
       .Y (n_1715));
  NAND4XL g180292(.A (n_1101), .B (n_1064), .C (n_1124), .D (n_1046),
       .Y (n_1714));
  AOI222X1 g180293(.A0 (n_970), .A1 (mem_rdata[22]), .B0
       (\reg_op1[6]_9643 ), .B1 (cpu_state[2]), .C0 (n_971), .C1
       (mem_rdata[14]), .Y (n_1713));
  NAND4XL g180294(.A (n_1128), .B (n_1131), .C (n_1105), .D (n_1130),
       .Y (n_1712));
  NAND4XL g180295(.A (n_1071), .B (n_1146), .C (n_1108), .D (n_1147),
       .Y (n_1711));
  NAND4XL g180296(.A (n_1040), .B (n_1126), .C (n_1053), .D (n_1039),
       .Y (n_1710));
  MX2X1 g180298(.A (\genblk1.pcpi_mul_rs1 [2]), .B (\reg_op1[2]_9639 ),
       .S0 (n_1310), .Y (n_1708));
  MX2X1 g180299(.A (\genblk1.pcpi_mul_rs1 [3]), .B (\reg_op1[3]_9640 ),
       .S0 (n_1310), .Y (n_1707));
  MX2X1 g180300(.A (\genblk1.pcpi_mul_rs1 [5]), .B (\reg_op1[5]_9642 ),
       .S0 (n_1310), .Y (n_1706));
  MX2X1 g180301(.A (\genblk1.pcpi_mul_rs1 [8]), .B (\reg_op1[8]_9645 ),
       .S0 (n_1310), .Y (n_1705));
  MX2X1 g180302(.A (\genblk1.pcpi_mul_rs1 [9]), .B (\reg_op1[9]_9646 ),
       .S0 (n_1310), .Y (n_1704));
  MX2X1 g180303(.A (\genblk1.pcpi_mul_rs1 [12]), .B (\reg_op1[12]_9649
       ), .S0 (n_1310), .Y (n_1703));
  MX2X1 g180304(.A (\genblk1.pcpi_mul_rs1 [14]), .B (\reg_op1[14]_9651
       ), .S0 (n_1310), .Y (n_1702));
  MX2X1 g180305(.A (\genblk1.pcpi_mul_rs1 [15]), .B (\reg_op1[15]_9652
       ), .S0 (n_1310), .Y (n_1701));
  MX2X1 g180306(.A (\genblk1.pcpi_mul_rs1 [10]), .B (\reg_op1[10]_9647
       ), .S0 (n_1310), .Y (n_1700));
  MX2X1 g180307(.A (\genblk1.pcpi_mul_rs1 [18]), .B (\reg_op1[18]_9655
       ), .S0 (n_1310), .Y (n_1699));
  MX2X1 g180308(.A (\genblk1.pcpi_mul_rs1 [19]), .B (\reg_op1[19]_9656
       ), .S0 (n_1310), .Y (n_1698));
  MX2X1 g180309(.A (\genblk1.pcpi_mul_rs1 [21]), .B (\reg_op1[21]_9658
       ), .S0 (n_1310), .Y (n_1697));
  MX2X1 g180310(.A (\genblk1.pcpi_mul_rs1 [22]), .B (\reg_op1[22]_9659
       ), .S0 (n_1310), .Y (n_1696));
  MX2X1 g180311(.A (\genblk1.pcpi_mul_rs1 [24]), .B (\reg_op1[24]_9661
       ), .S0 (n_1310), .Y (n_1695));
  MX2X1 g180312(.A (\genblk1.pcpi_mul_rs1 [25]), .B (\reg_op1[25]_9662
       ), .S0 (n_1310), .Y (n_1694));
  MX2X1 g180313(.A (\genblk1.pcpi_mul_rs1 [27]), .B (\reg_op1[27]_9664
       ), .S0 (n_1310), .Y (n_1693));
  MX2X1 g180314(.A (\genblk1.pcpi_mul_rs1 [30]), .B (\reg_op1[30]_9667
       ), .S0 (n_1310), .Y (n_1692));
  MX2X1 g180315(.A (\genblk1.pcpi_mul_rs1 [1]), .B (\reg_op1[1]_9638 ),
       .S0 (n_1310), .Y (n_1691));
  MX2X1 g180316(.A (\genblk1.pcpi_mul_rs2 [4]), .B (\reg_op2[4]_9673 ),
       .S0 (n_1310), .Y (n_1690));
  MX2X1 g180317(.A (\genblk1.pcpi_mul_rs2 [14]), .B (\reg_op2[14]_9683
       ), .S0 (n_1310), .Y (n_1689));
  MX2X1 g180318(.A (\genblk1.pcpi_mul_rs2 [16]), .B (\reg_op2[16]_9685
       ), .S0 (n_1310), .Y (n_1688));
  MX2X1 g180319(.A (\genblk1.pcpi_mul_rs2 [18]), .B (\reg_op2[18]_9687
       ), .S0 (n_1310), .Y (n_1687));
  MX2X1 g180320(.A (\genblk1.pcpi_mul_rs2 [20]), .B (\reg_op2[20]_9689
       ), .S0 (n_1310), .Y (n_1686));
  MX2X1 g180321(.A (\genblk1.pcpi_mul_rs2 [22]), .B (\reg_op2[22]_9691
       ), .S0 (n_1310), .Y (n_1685));
  MX2X1 g180322(.A (\genblk1.pcpi_mul_rs2 [24]), .B (\reg_op2[24]_9693
       ), .S0 (n_1310), .Y (n_1684));
  MX2X1 g180323(.A (\genblk1.pcpi_mul_rs2 [26]), .B (\reg_op2[26]_9695
       ), .S0 (n_1310), .Y (n_1683));
  MX2X1 g180324(.A (\genblk1.pcpi_mul_rs2 [28]), .B (\reg_op2[28]_9697
       ), .S0 (n_1310), .Y (n_1682));
  MX2X1 g180325(.A (\genblk1.pcpi_mul_rs2 [30]), .B (\reg_op2[30]_9699
       ), .S0 (n_1310), .Y (n_1681));
  MX2X1 g180326(.A (\genblk1.pcpi_mul_rs2 [6]), .B (\reg_op2[6]_9675 ),
       .S0 (n_1310), .Y (n_1680));
  MX2X1 g180327(.A (\genblk1.pcpi_mul_rs2 [0]), .B (\reg_op2[0]_9669 ),
       .S0 (n_1310), .Y (n_1679));
  MX2X1 g180328(.A (\genblk1.pcpi_mul_rs1 [23]), .B (\reg_op1[23]_9660
       ), .S0 (n_1310), .Y (n_1678));
  MX2X1 g180329(.A (\genblk1.pcpi_mul_rs1 [6]), .B (\reg_op1[6]_9643 ),
       .S0 (n_1310), .Y (n_1677));
  MX2X1 g180330(.A (\genblk1.pcpi_mul_rs1 [13]), .B (\reg_op1[13]_9650
       ), .S0 (n_1310), .Y (n_1676));
  MX2X1 g180331(.A (\genblk1.pcpi_mul_rs1 [26]), .B (\reg_op1[26]_9663
       ), .S0 (n_1310), .Y (n_1675));
  MX2X1 g180332(.A (\genblk1.pcpi_mul_rs2 [12]), .B (\reg_op2[12]_9681
       ), .S0 (n_1310), .Y (n_1674));
  MX2X1 g180333(.A (\genblk1.pcpi_mul_rs2 [10]), .B (\reg_op2[10]_9679
       ), .S0 (n_1310), .Y (n_1673));
  MX2X1 g180334(.A (\genblk1.pcpi_mul_rs1 [7]), .B (\reg_op1[7]_9644 ),
       .S0 (n_1310), .Y (n_1672));
  MX2X1 g180335(.A (\genblk1.pcpi_mul_rs2 [8]), .B (\reg_op2[8]_9677 ),
       .S0 (n_1310), .Y (n_1671));
  MX2X1 g180336(.A (\genblk1.pcpi_mul_rs1 [11]), .B (\reg_op1[11]_9648
       ), .S0 (n_1310), .Y (n_1670));
  MX2X1 g180337(.A (\genblk1.pcpi_mul_rs1 [4]), .B (\reg_op1[4]_9641 ),
       .S0 (n_1310), .Y (n_1669));
  MX2X1 g180338(.A (\genblk1.pcpi_mul_rs1 [16]), .B (\reg_op1[16]_9653
       ), .S0 (n_1310), .Y (n_1668));
  MX2X1 g180339(.A (\genblk1.pcpi_mul_rs1 [20]), .B (\reg_op1[20]_9657
       ), .S0 (n_1310), .Y (n_1667));
  MX2X1 g180340(.A (\genblk1.pcpi_mul_rs1 [28]), .B (\reg_op1[28]_9665
       ), .S0 (n_1310), .Y (n_1666));
  MX2X1 g180341(.A (\genblk1.pcpi_mul_rs1 [29]), .B (\reg_op1[29]_9666
       ), .S0 (n_1310), .Y (n_1665));
  MX2X1 g180342(.A (\genblk1.pcpi_mul_rs2 [2]), .B (\reg_op2[2]_9671 ),
       .S0 (n_1310), .Y (n_1664));
  MX2X1 g180343(.A (\genblk1.pcpi_mul_rs1 [31]), .B (\reg_op1[31]_9668
       ), .S0 (n_1310), .Y (n_1663));
  MX2X1 g180344(.A (\genblk1.pcpi_mul_rs1 [17]), .B (\reg_op1[17]_9654
       ), .S0 (n_1310), .Y (n_1662));
  MX2X1 g180345(.A (\reg_op2[0]_9669 ), .B (n_5630), .S0 (n_542), .Y
       (n_1661));
  MX2X1 g180346(.A (\reg_op2[1]_9670 ), .B (n_5631), .S0 (n_542), .Y
       (n_1660));
  MX2X1 g180347(.A (\reg_op2[2]_9671 ), .B (n_5632), .S0 (n_542), .Y
       (n_1659));
  MX2X1 g180348(.A (\reg_op2[3]_9672 ), .B (n_5633), .S0 (n_542), .Y
       (n_1658));
  MX2X1 g180349(.A (\reg_op2[4]_9673 ), .B (n_5634), .S0 (n_542), .Y
       (n_1657));
  MX2X1 g180350(.A (\reg_op2[5]_9674 ), .B (n_5635), .S0 (n_542), .Y
       (n_1656));
  MX2X1 g180351(.A (\reg_op2[6]_9675 ), .B (n_5636), .S0 (n_542), .Y
       (n_1655));
  MX2X1 g180352(.A (\reg_op2[7]_9676 ), .B (n_5637), .S0 (n_542), .Y
       (n_1654));
  AOI222X1 g180366(.A0 (mem_rdata_q[10]), .A1 (n_505), .B0
       (mem_rdata[10]), .B1 (n_839), .C0 (n_562), .C1 (n_1203), .Y
       (n_1816));
  MX2X1 g180367(.A (n_1214), .B (n_1362), .S0 (mem_la_secondword), .Y
       (n_1815));
  OAI2BB1X1 g180368(.A0N (n_562), .A1N (n_1207), .B0 (n_1431), .Y
       (n_1814));
  OAI221X1 g180369(.A0 (mem_la_secondword), .A1 (n_1213), .B0 (n_643),
       .B1 (n_663), .C0 (n_1271), .Y (n_1813));
  OAI221X1 g180370(.A0 (mem_la_secondword), .A1 (n_1211), .B0 (n_649),
       .B1 (n_663), .C0 (n_1281), .Y (n_1812));
  OAI221X1 g180371(.A0 (mem_la_secondword), .A1 (n_1202), .B0 (n_594),
       .B1 (n_663), .C0 (n_1234), .Y (n_1811));
  OAI221X1 g180372(.A0 (mem_la_secondword), .A1 (n_1206), .B0 (n_586),
       .B1 (n_663), .C0 (n_1256), .Y (n_1810));
  AOI221X1 g180373(.A0 (mem_rdata_q[15]), .A1 (n_505), .B0
       (mem_rdata[15]), .B1 (n_839), .C0 (n_1533), .Y (n_1809));
  AOI222X1 g180374(.A0 (mem_rdata_q[11]), .A1 (n_505), .B0
       (mem_rdata[11]), .B1 (n_839), .C0 (n_562), .C1 (n_1205), .Y
       (n_1808));
  AOI221X1 g180375(.A0 (mem_rdata_q[8]), .A1 (n_505), .B0
       (mem_rdata[8]), .B1 (n_839), .C0 (n_1528), .Y (n_1807));
  MX2X1 g180376(.A (n_1208), .B (n_1197), .S0 (mem_la_secondword), .Y
       (n_1806));
  OAI22X1 g180377(.A0 (mem_la_secondword), .A1 (n_1201), .B0 (n_562),
       .B1 (n_1204), .Y (n_1805));
  AOI221X1 g180378(.A0 (mem_rdata_q[9]), .A1 (n_505), .B0
       (mem_rdata[9]), .B1 (n_839), .C0 (n_1544), .Y (n_1804));
  AOI221X1 g180379(.A0 (mem_rdata_q[2]), .A1 (n_505), .B0
       (mem_rdata[2]), .B1 (n_839), .C0 (n_1526), .Y (n_1803));
  AOI222X1 g180380(.A0 (mem_rdata[0]), .A1 (n_839), .B0
       (mem_rdata_q[0]), .B1 (n_505), .C0 (n_562), .C1 (n_6864), .Y
       (n_1802));
  INVX1 g180381(.A (n_1623), .Y (n_1624));
  INVX1 g180384(.A (n_1617), .Y (n_1618));
  INVX1 g180385(.A (n_1615), .Y (n_1616));
  INVX1 g180386(.A (n_11745), .Y (n_1613));
  INVX1 g180387(.A (n_1609), .Y (n_1610));
  INVX1 g180389(.A (n_1600), .Y (n_1601));
  INVX1 g180390(.A (n_1590), .Y (n_1589));
  INVX1 g180391(.A (n_1585), .Y (n_1584));
  AOI222X1 g180412(.A0 (count_cycle[33]), .A1 (instr_rdcycleh), .B0
       (count_cycle[1]), .B1 (instr_rdcycle), .C0
       (\genblk1.pcpi_mul_rd [33]), .C1 (n_11690), .Y (n_1560));
  NOR4X1 g180413(.A (n_6673), .B (n_6659), .C (n_6657), .D (n_1165), .Y
       (n_1559));
  OAI2BB1X1 g180414(.A0N (instr_sb), .A1N (cpu_state[1]), .B0 (n_1306),
       .Y (n_1558));
  OAI2BB1X1 g180415(.A0N (instr_sh), .A1N (cpu_state[1]), .B0 (n_1272),
       .Y (n_1557));
  NAND3BXL g180416(.AN (n_5597), .B (n_5598), .C (n_1310), .Y (n_1556));
  OAI2BB1X1 g180417(.A0N (compressed_instr), .A1N (n_953), .B0 (n_335),
       .Y (n_1555));
  NAND3X1 g180418(.A (decoded_rd[4]), .B (cpu_state[6]), .C (n_1319),
       .Y (n_1554));
  OAI2BB1X1 g180419(.A0N (pcpi_timeout_counter[3]), .A1N (n_218), .B0
       (n_307), .Y (n_1553));
  NAND3X1 g180420(.A (decoded_rd[0]), .B (cpu_state[6]), .C (n_1319),
       .Y (n_1552));
  NOR2X1 g180422(.A (n_1166), .B (n_544), .Y (n_1550));
  NAND2X1 g180423(.A (n_613), .B (n_1355), .Y (n_1549));
  NAND2X1 g180424(.A (n_279), .B (n_1347), .Y (n_1548));
  NAND2X1 g180425(.A (n_279), .B (n_1348), .Y (n_1547));
  NAND2X1 g180426(.A (n_279), .B (n_1354), .Y (n_1546));
  NAND2X1 g180427(.A (n_279), .B (n_1346), .Y (n_1545));
  NOR2X1 g180428(.A (mem_la_secondword), .B (n_1210), .Y (n_1544));
  NAND2X1 g180429(.A (latched_is_lh), .B (n_1199), .Y (n_1543));
  NAND2X1 g180430(.A (n_279), .B (n_1353), .Y (n_1542));
  OAI2BB1X1 g180431(.A0N (n_871), .A1N (n_6548), .B0 (n_136), .Y
       (n_1541));
  OAI2BB1X1 g180432(.A0N (n_770), .A1N (n_258), .B0 (n_307), .Y
       (n_1540));
  NAND2X1 g180433(.A (decoded_imm[24]), .B (n_421), .Y (n_1539));
  NAND2X1 g180434(.A (decoded_imm[7]), .B (n_421), .Y (n_1538));
  NAND2X1 g180435(.A (mem_rdata_q[11]), .B (n_1328), .Y (n_1537));
  NOR2BX1 g180436(.AN (alu_out_q[0]), .B (n_11742), .Y (n_1536));
  NAND2X1 g180437(.A (n_985), .B (n_1339), .Y (n_1535));
  OR2X1 g180438(.A (mem_rdata_q[16]), .B (n_1215), .Y (n_1534));
  NOR2X1 g180439(.A (mem_la_secondword), .B (n_1200), .Y (n_1533));
  NAND2X1 g180440(.A (mem_rdata_q[10]), .B (n_1328), .Y (n_1532));
  NAND2X1 g180441(.A (reg_pc[23]), .B (n_547), .Y (n_1531));
  NAND2X1 g180442(.A (n_2), .B (n_52), .Y (n_1530));
  NOR2BX1 g180443(.AN (n_993), .B (n_676), .Y (n_1529));
  NOR2X1 g180444(.A (mem_la_secondword), .B (n_1212), .Y (n_1528));
  NAND2X1 g180445(.A (decoded_imm[29]), .B (n_421), .Y (n_1527));
  NOR2X1 g180446(.A (mem_la_secondword), .B (n_1209), .Y (n_1526));
  NOR2X1 g180447(.A (reg_sh[2]), .B (n_1322), .Y (n_1525));
  NAND2X1 g180456(.A (n_676), .B (n_1340), .Y (n_1640));
  NAND2X1 g180461(.A (n_983), .B (n_1343), .Y (n_1639));
  NOR2X1 g180464(.A (n_356), .B (n_1339), .Y (n_1638));
  NAND3BXL g180476(.AN (n_5598), .B (n_5597), .C (n_1310), .Y (n_1637));
  NAND3BXL g180479(.AN (n_881), .B (cpu_state[0]), .C (n_582), .Y
       (n_1636));
  NAND3BXL g180482(.AN (n_986), .B (n_6542), .C (n_152), .Y (n_1635));
  OR2X1 g180484(.A (n_1321), .B (n_1325), .Y (n_1634));
  AND3XL g180485(.A (n_599), .B (n_981), .C (n_973), .Y (n_1633));
  NAND2BX1 g180488(.AN (n_1193), .B (n_1369), .Y (n_1632));
  NOR2X1 g180489(.A (n_611), .B (n_1322), .Y (n_1631));
  NAND2X1 g180490(.A (n_545), .B (n_1193), .Y (n_1630));
  NOR2X1 g180491(.A (reg_sh[0]), .B (n_676), .Y (n_1629));
  OR2X1 g180492(.A (mem_do_wdata), .B (n_1341), .Y (n_1628));
  NOR2X1 g180497(.A (n_289), .B (n_1332), .Y (n_1627));
  NOR2X1 g180498(.A (n_963), .B (n_1334), .Y (n_1626));
  NOR2X1 g180499(.A (n_289), .B (n_1334), .Y (n_1625));
  NAND2X1 g180500(.A (n_962), .B (n_1333), .Y (n_1623));
  NOR2BX1 g180501(.AN (n_1333), .B (n_338), .Y (n_1622));
  AND2X1 g180502(.A (n_1335), .B (n_962), .Y (n_1621));
  NOR2BX1 g180503(.AN (n_1364), .B (mem_rdata_latched[0]), .Y (n_1620));
  NOR2X1 g180504(.A (n_974), .B (n_335), .Y (n_1619));
  NAND2X1 g180505(.A (n_962), .B (n_8), .Y (n_1617));
  NAND2X1 g180507(.A (n_665), .B (n_8), .Y (n_1615));
  NOR2X1 g180508(.A (n_289), .B (n_1336), .Y (n_1614));
  NOR2X1 g180511(.A (n_963), .B (n_1336), .Y (n_1611));
  NAND2X1 g180512(.A (n_842), .B (n_8), .Y (n_1609));
  NOR2X1 g180513(.A (n_843), .B (n_7), .Y (n_1608));
  NOR2X1 g180515(.A (n_963), .B (n_7), .Y (n_1607));
  NOR2X1 g180516(.A (n_843), .B (n_1336), .Y (n_1606));
  NOR2X1 g180517(.A (n_289), .B (n_7), .Y (n_1605));
  NOR2X1 g180519(.A (n_338), .B (n_1345), .Y (n_1604));
  AND2X1 g180520(.A (n_1333), .B (n_665), .Y (n_1603));
  NOR2X1 g180521(.A (n_963), .B (n_1332), .Y (n_1602));
  NAND2X1 g180522(.A (n_842), .B (n_1335), .Y (n_1600));
  NOR2X1 g180523(.A (n_338), .B (n_1336), .Y (n_1599));
  NOR2X1 g180524(.A (n_338), .B (n_7), .Y (n_1598));
  AND2X1 g180525(.A (n_1333), .B (n_842), .Y (n_1597));
  NOR2X1 g180526(.A (n_289), .B (n_1345), .Y (n_1596));
  NOR2X1 g180527(.A (n_843), .B (n_1345), .Y (n_1595));
  NOR2X1 g180528(.A (n_338), .B (n_1334), .Y (n_1594));
  NOR2X1 g180529(.A (n_843), .B (n_1332), .Y (n_1593));
  NOR2X1 g180530(.A (n_338), .B (n_1332), .Y (n_1592));
  NOR2X1 g180531(.A (n_843), .B (n_1334), .Y (n_1591));
  NAND2X1 g180533(.A (mem_rdata_latched[0]), .B (n_1364), .Y (n_1590));
  NOR2X1 g180534(.A (n_345), .B (n_335), .Y (n_1588));
  AND2X2 g180535(.A (n_1368), .B (n_668), .Y (n_434));
  OR2X2 g180536(.A (n_427), .B (n_1191), .Y (n_1586));
  OR2X1 g180537(.A (n_1368), .B (n_954), .Y (n_1585));
  AO22X2 g180538(.A0 (n_442), .A1 (n_208), .B0 (latched_branch), .B1
       (n_6704), .Y (n_406));
  AND2X2 g180539(.A (n_1367), .B (n_668), .Y (n_460));
  AND2X2 g180540(.A (n_542), .B (n_1370), .Y (n_472));
  INVX2 g180541(.A (n_1517), .Y (n_1518));
  INVX2 g180542(.A (n_1514), .Y (n_1515));
  INVX2 g180543(.A (n_1512), .Y (n_1513));
  AOI22X1 g180544(.A0 (decoded_imm_j[4]), .A1 (n_441), .B0
       (decoded_imm[4]), .B1 (n_537), .Y (n_1488));
  MX2X1 g180550(.A (compressed_instr), .B (latched_compr), .S0 (n_324),
       .Y (n_1482));
  AOI22XL g180552(.A0 (n_666), .A1 (n_7026), .B0 (count_instr[29]), .B1
       (n_952), .Y (n_1480));
  AOI22XL g180553(.A0 (n_666), .A1 (n_7047), .B0 (count_instr[8]), .B1
       (n_952), .Y (n_1479));
  AOI22XL g180554(.A0 (n_666), .A1 (n_7049), .B0 (count_instr[6]), .B1
       (n_952), .Y (n_1478));
  AOI22XL g180555(.A0 (n_666), .A1 (n_7030), .B0 (count_instr[25]), .B1
       (n_952), .Y (n_1477));
  AOI22X1 g180556(.A0 (decoded_imm_j[3]), .A1 (n_441), .B0
       (decoded_imm[3]), .B1 (n_537), .Y (n_1476));
  AOI22XL g180557(.A0 (n_666), .A1 (n_7034), .B0 (count_instr[21]), .B1
       (n_952), .Y (n_1475));
  AOI22XL g180558(.A0 (n_666), .A1 (n_7036), .B0 (count_instr[19]), .B1
       (n_952), .Y (n_1474));
  AOI22XL g180559(.A0 (n_666), .A1 (n_7037), .B0 (count_instr[18]), .B1
       (n_952), .Y (n_1473));
  AOI22XL g180560(.A0 (n_666), .A1 (n_7018), .B0 (count_instr[37]), .B1
       (n_952), .Y (n_1472));
  AOI22XL g180562(.A0 (n_666), .A1 (n_7017), .B0 (count_instr[38]), .B1
       (n_952), .Y (n_1470));
  AOI22XL g180563(.A0 (n_666), .A1 (n_7016), .B0 (count_instr[39]), .B1
       (n_952), .Y (n_1469));
  AOI22XL g180564(.A0 (n_666), .A1 (n_7015), .B0 (count_instr[40]), .B1
       (n_952), .Y (n_1468));
  AOI22X1 g180565(.A0 (n_833), .A1 (n_52), .B0 (reg_pc[30]), .B1
       (n_961), .Y (n_1467));
  AOI22XL g180566(.A0 (n_666), .A1 (n_7052), .B0 (count_instr[3]), .B1
       (n_952), .Y (n_1466));
  AOI22X1 g180567(.A0 (decoded_imm_j[12]), .A1 (n_441), .B0
       (decoded_imm[12]), .B1 (n_537), .Y (n_1465));
  AOI22X1 g180568(.A0 (decoded_imm_j[1]), .A1 (n_441), .B0
       (decoded_imm[1]), .B1 (n_537), .Y (n_1464));
  AOI22X1 g180570(.A0 (decoded_imm_j[8]), .A1 (n_441), .B0
       (decoded_imm[8]), .B1 (n_537), .Y (n_1462));
  AOI22XL g180571(.A0 (n_666), .A1 (n_7012), .B0 (count_instr[43]), .B1
       (n_952), .Y (n_1461));
  AOI22X1 g180572(.A0 (decoded_imm_j[2]), .A1 (n_441), .B0
       (decoded_imm[2]), .B1 (n_537), .Y (n_1460));
  AOI22X1 g180573(.A0 (n_833), .A1 (n_64), .B0 (reg_pc[2]), .B1
       (n_961), .Y (n_1459));
  AO22X1 g180574(.A0 (n_833), .A1 (n_114), .B0 (reg_pc[3]), .B1
       (n_961), .Y (n_1458));
  AOI22XL g180575(.A0 (n_666), .A1 (n_7011), .B0 (count_instr[44]), .B1
       (n_952), .Y (n_1457));
  AOI22XL g180576(.A0 (n_972), .A1 (mem_rdata[2]), .B0 (cpu_state[3]),
       .B1 (n_6990), .Y (n_1456));
  AOI22X1 g180577(.A0 (decoded_imm_j[13]), .A1 (n_441), .B0
       (decoded_imm[13]), .B1 (n_537), .Y (n_1455));
  AOI22XL g180578(.A0 (n_972), .A1 (mem_rdata[5]), .B0 (cpu_state[3]),
       .B1 (n_6987), .Y (n_1454));
  AOI22XL g180579(.A0 (n_666), .A1 (n_7014), .B0 (count_instr[41]), .B1
       (n_952), .Y (n_1453));
  AOI22XL g180580(.A0 (n_666), .A1 (n_7043), .B0 (count_instr[12]), .B1
       (n_952), .Y (n_1452));
  AOI22XL g180581(.A0 (n_666), .A1 (n_7025), .B0 (count_instr[30]), .B1
       (n_952), .Y (n_1451));
  AOI22XL g180583(.A0 (n_666), .A1 (n_7005), .B0 (count_instr[50]), .B1
       (n_952), .Y (n_1449));
  AOI22X1 g180584(.A0 (n_833), .A1 (n_68), .B0 (reg_pc[31]), .B1
       (n_961), .Y (n_1448));
  AOI22XL g180585(.A0 (n_972), .A1 (mem_rdata[3]), .B0 (cpu_state[3]),
       .B1 (n_6989), .Y (n_1447));
  AOI22XL g180586(.A0 (n_972), .A1 (mem_rdata[6]), .B0 (cpu_state[3]),
       .B1 (n_6986), .Y (n_1446));
  AOI22X1 g180587(.A0 (decoded_imm_j[17]), .A1 (n_441), .B0
       (decoded_imm[17]), .B1 (n_537), .Y (n_1445));
  AOI22XL g180588(.A0 (n_666), .A1 (n_7053), .B0 (count_instr[2]), .B1
       (n_952), .Y (n_1444));
  AOI22X1 g180589(.A0 (decoded_imm_j[11]), .A1 (n_441), .B0
       (decoded_imm[11]), .B1 (n_537), .Y (n_1443));
  AOI22X1 g180590(.A0 (decoded_imm_j[14]), .A1 (n_441), .B0
       (decoded_imm[14]), .B1 (n_537), .Y (n_1442));
  AOI22XL g180591(.A0 (n_666), .A1 (n_7013), .B0 (count_instr[42]), .B1
       (n_952), .Y (n_1441));
  AOI22XL g180592(.A0 (n_666), .A1 (n_7051), .B0 (count_instr[4]), .B1
       (n_952), .Y (n_1440));
  AOI22XL g180594(.A0 (n_972), .A1 (mem_rdata[4]), .B0 (cpu_state[3]),
       .B1 (n_6988), .Y (n_1438));
  AOI22XL g180595(.A0 (n_666), .A1 (n_7054), .B0 (count_instr[1]), .B1
       (n_952), .Y (n_1437));
  AOI22XL g180596(.A0 (n_666), .A1 (n_7040), .B0 (count_instr[15]), .B1
       (n_952), .Y (n_1436));
  AOI22XL g180597(.A0 (n_666), .A1 (n_7050), .B0 (count_instr[5]), .B1
       (n_952), .Y (n_1435));
  AOI22XL g180598(.A0 (n_666), .A1 (n_7041), .B0 (count_instr[14]), .B1
       (n_952), .Y (n_1434));
  AOI22X1 g180599(.A0 (decoded_imm_j[9]), .A1 (n_441), .B0
       (decoded_imm[9]), .B1 (n_537), .Y (n_1433));
  AOI22XL g180600(.A0 (n_666), .A1 (n_7031), .B0 (count_instr[24]), .B1
       (n_952), .Y (n_1432));
  AOI22X1 g180601(.A0 (mem_rdata_q[12]), .A1 (n_505), .B0
       (mem_rdata[12]), .B1 (n_839), .Y (n_1431));
  AOI22XL g180602(.A0 (n_666), .A1 (n_7035), .B0 (count_instr[20]), .B1
       (n_952), .Y (n_1430));
  AOI22X1 g180604(.A0 (decoded_imm_j[15]), .A1 (n_441), .B0
       (decoded_imm[15]), .B1 (n_537), .Y (n_1428));
  AOI22X1 g180605(.A0 (decoded_imm_j[16]), .A1 (n_441), .B0
       (decoded_imm[16]), .B1 (n_537), .Y (n_1427));
  AOI22X1 g180606(.A0 (decoded_imm_j[18]), .A1 (n_441), .B0
       (decoded_imm[18]), .B1 (n_537), .Y (n_1426));
  AOI22X1 g180607(.A0 (decoded_imm_j[19]), .A1 (n_441), .B0
       (decoded_imm[19]), .B1 (n_537), .Y (n_1425));
  AOI22XL g180608(.A0 (n_666), .A1 (n_7033), .B0 (count_instr[22]), .B1
       (n_952), .Y (n_1424));
  OAI211X1 g180609(.A0 (\reg_op1[27]_9664 ), .A1 (n_760), .B0
       (\reg_op1[26]_9663 ), .C0 (\genblk2.pcpi_div_minus_2470_59_n_488
       ), .Y (n_1423));
  AOI32X1 g180610(.A0 (\reg_op1[24]_9661 ), .A1
       (\genblk2.pcpi_div_minus_2470_59_n_483 ), .A2 (n_156), .B0
       (\reg_op1[25]_9662 ), .B1 (n_722), .Y (n_1422));
  AOI32X1 g180611(.A0 (\reg_op1[16]_9653 ), .A1
       (\genblk2.pcpi_div_minus_2470_59_n_481 ), .A2 (n_154), .B0
       (\reg_op1[17]_9654 ), .B1 (n_726), .Y (n_1421));
  XNOR2X1 g180612(.A (count_instr[0]), .B (n_666), .Y (n_1420));
  AOI32X1 g180613(.A0 (\reg_op2[14]_9683 ), .A1 (\reg_op1[14]_9651 ),
       .A2 (n_283), .B0 (is_lui_auipc_jal_jalr_addi_add_sub), .B1
       (n_6639), .Y (n_1419));
  NOR4X1 g180614(.A (\reg_op2[21]_9690 ), .B (\reg_op2[3]_9672 ), .C
       (\reg_op2[22]_9691 ), .D (\reg_op2[23]_9692 ), .Y (n_1418));
  AOI32X1 g180615(.A0 (\reg_op2[18]_9687 ), .A1 (\reg_op1[18]_9655 ),
       .A2 (n_283), .B0 (is_lui_auipc_jal_jalr_addi_add_sub), .B1
       (n_6643), .Y (n_1417));
  AOI32X1 g180616(.A0 (\reg_op2[8]_9677 ), .A1 (\reg_op1[8]_9645 ), .A2
       (n_283), .B0 (is_lui_auipc_jal_jalr_addi_add_sub), .B1 (n_6633),
       .Y (n_1416));
  AOI32X1 g180617(.A0 (\reg_op2[7]_9676 ), .A1 (\reg_op1[7]_9644 ), .A2
       (n_283), .B0 (is_lui_auipc_jal_jalr_addi_add_sub), .B1 (n_6632),
       .Y (n_1415));
  AOI32X1 g180618(.A0 (\reg_op2[6]_9675 ), .A1 (\reg_op1[6]_9643 ), .A2
       (n_283), .B0 (is_lui_auipc_jal_jalr_addi_add_sub), .B1 (n_6631),
       .Y (n_1414));
  AOI32X1 g180619(.A0 (\reg_op2[10]_9679 ), .A1 (\reg_op1[10]_9647 ),
       .A2 (n_283), .B0 (is_lui_auipc_jal_jalr_addi_add_sub), .B1
       (n_6635), .Y (n_1413));
  AOI22XL g180620(.A0 (n_666), .A1 (n_6997), .B0 (count_instr[58]), .B1
       (n_952), .Y (n_1412));
  AOI221X1 g180621(.A0 (n_607), .A1 (mem_rdata[1]), .B0 (n_340), .B1
       (mem_rdata[17]), .C0 (n_1125), .Y (n_1411));
  AOI32X1 g180622(.A0 (\reg_op2[13]_9682 ), .A1 (\reg_op1[13]_9650 ),
       .A2 (n_283), .B0 (is_lui_auipc_jal_jalr_addi_add_sub), .B1
       (n_6638), .Y (n_1410));
  AOI32X1 g180623(.A0 (\reg_op2[11]_9680 ), .A1 (\reg_op1[11]_9648 ),
       .A2 (n_283), .B0 (is_lui_auipc_jal_jalr_addi_add_sub), .B1
       (n_6636), .Y (n_1409));
  AOI32X1 g180624(.A0 (\reg_op2[9]_9678 ), .A1 (\reg_op1[9]_9646 ), .A2
       (n_283), .B0 (is_lui_auipc_jal_jalr_addi_add_sub), .B1 (n_6634),
       .Y (n_1408));
  AOI32X1 g180625(.A0 (\reg_op2[15]_9684 ), .A1 (\reg_op1[15]_9652 ),
       .A2 (n_283), .B0 (is_lui_auipc_jal_jalr_addi_add_sub), .B1
       (n_6640), .Y (n_1407));
  AOI32X1 g180626(.A0 (\reg_op2[12]_9681 ), .A1 (\reg_op1[12]_9649 ),
       .A2 (n_283), .B0 (is_lui_auipc_jal_jalr_addi_add_sub), .B1
       (n_6637), .Y (n_1406));
  AOI22XL g180627(.A0 (n_666), .A1 (n_7021), .B0 (count_instr[34]), .B1
       (n_952), .Y (n_1405));
  AOI22XL g180628(.A0 (n_666), .A1 (n_7022), .B0 (count_instr[33]), .B1
       (n_952), .Y (n_1404));
  AOI22XL g180629(.A0 (n_666), .A1 (n_7010), .B0 (count_instr[45]), .B1
       (n_952), .Y (n_1403));
  AOI22XL g180630(.A0 (n_666), .A1 (n_7009), .B0 (count_instr[46]), .B1
       (n_952), .Y (n_1402));
  AOI22XL g180631(.A0 (n_666), .A1 (n_7008), .B0 (count_instr[47]), .B1
       (n_952), .Y (n_1401));
  AOI22XL g180632(.A0 (n_666), .A1 (n_7007), .B0 (count_instr[48]), .B1
       (n_952), .Y (n_1400));
  AOI22XL g180633(.A0 (n_666), .A1 (n_7006), .B0 (count_instr[49]), .B1
       (n_952), .Y (n_1399));
  AOI22XL g180634(.A0 (n_666), .A1 (n_7004), .B0 (count_instr[51]), .B1
       (n_952), .Y (n_1398));
  AOI22XL g180635(.A0 (n_666), .A1 (n_7003), .B0 (count_instr[52]), .B1
       (n_952), .Y (n_1397));
  AOI22XL g180636(.A0 (n_666), .A1 (n_7001), .B0 (count_instr[54]), .B1
       (n_952), .Y (n_1396));
  AOI22XL g180637(.A0 (n_666), .A1 (n_7002), .B0 (count_instr[53]), .B1
       (n_952), .Y (n_1395));
  AOI22XL g180638(.A0 (n_666), .A1 (n_6999), .B0 (count_instr[56]), .B1
       (n_952), .Y (n_1394));
  AOI22XL g180639(.A0 (n_666), .A1 (n_6998), .B0 (count_instr[57]), .B1
       (n_952), .Y (n_1393));
  AOI22XL g180640(.A0 (n_666), .A1 (n_6996), .B0 (count_instr[59]), .B1
       (n_952), .Y (n_1392));
  AOI22XL g180641(.A0 (n_666), .A1 (n_6995), .B0 (count_instr[60]), .B1
       (n_952), .Y (n_1391));
  AOI22XL g180642(.A0 (n_666), .A1 (n_6994), .B0 (count_instr[61]), .B1
       (n_952), .Y (n_1390));
  AOI22XL g180643(.A0 (n_666), .A1 (n_6993), .B0 (count_instr[62]), .B1
       (n_952), .Y (n_1389));
  AOI22XL g180644(.A0 (n_666), .A1 (n_7023), .B0 (count_instr[32]), .B1
       (n_952), .Y (n_1388));
  AOI22XL g180645(.A0 (n_666), .A1 (n_6992), .B0 (count_instr[63]), .B1
       (n_952), .Y (n_1387));
  AOI22XL g180646(.A0 (n_666), .A1 (n_7028), .B0 (count_instr[27]), .B1
       (n_952), .Y (n_1386));
  AOI22XL g180647(.A0 (n_666), .A1 (n_7020), .B0 (count_instr[35]), .B1
       (n_952), .Y (n_1385));
  AOI22XL g180648(.A0 (n_666), .A1 (n_7048), .B0 (count_instr[7]), .B1
       (n_952), .Y (n_1384));
  AOI22XL g180649(.A0 (n_666), .A1 (n_7024), .B0 (count_instr[31]), .B1
       (n_952), .Y (n_1383));
  AOI22XL g180650(.A0 (n_666), .A1 (n_7000), .B0 (count_instr[55]), .B1
       (n_952), .Y (n_1382));
  AOI22XL g180651(.A0 (n_666), .A1 (n_7044), .B0 (count_instr[11]), .B1
       (n_952), .Y (n_1381));
  AOI22XL g180652(.A0 (n_666), .A1 (n_7019), .B0 (count_instr[36]), .B1
       (n_952), .Y (n_1380));
  AOI22XL g180653(.A0 (n_666), .A1 (n_7039), .B0 (count_instr[16]), .B1
       (n_952), .Y (n_1379));
  AOI22XL g180654(.A0 (n_666), .A1 (n_7027), .B0 (count_instr[28]), .B1
       (n_952), .Y (n_1378));
  AOI22XL g180655(.A0 (n_666), .A1 (n_7029), .B0 (count_instr[26]), .B1
       (n_952), .Y (n_1377));
  AOI22XL g180656(.A0 (n_666), .A1 (n_7042), .B0 (count_instr[13]), .B1
       (n_952), .Y (n_1376));
  AOI22XL g180657(.A0 (n_666), .A1 (n_7045), .B0 (count_instr[10]), .B1
       (n_952), .Y (n_1375));
  AOI22XL g180658(.A0 (n_666), .A1 (n_7038), .B0 (count_instr[17]), .B1
       (n_952), .Y (n_1374));
  AOI22XL g180659(.A0 (n_666), .A1 (n_7032), .B0 (count_instr[23]), .B1
       (n_952), .Y (n_1373));
  AOI22XL g180660(.A0 (n_666), .A1 (n_7046), .B0 (count_instr[9]), .B1
       (n_952), .Y (n_1372));
  AOI221X1 g180661(.A0 (n_657), .A1 (mem_rdata[15]), .B0 (n_340), .B1
       (mem_rdata[23]), .C0 (n_1094), .Y (n_1523));
  NOR4X1 g180662(.A (instr_rdinstrh), .B (instr_rdinstr), .C
       (instr_rdcycle), .D (instr_rdcycleh), .Y (n_288));
  AO22X2 g180663(.A0 (n_442), .A1 (n_160), .B0 (latched_branch), .B1
       (n_6678), .Y (n_398));
  AO22X2 g180664(.A0 (n_442), .A1 (n_164), .B0 (latched_branch), .B1
       (n_6682), .Y (n_394));
  AO22X2 g180665(.A0 (n_442), .A1 (n_196), .B0 (latched_branch), .B1
       (n_6695), .Y (n_382));
  AOI22XL g180666(.A0 (n_442), .A1 (n_142), .B0 (latched_branch), .B1
       (n_6696), .Y (n_1517));
  AO22X2 g180667(.A0 (n_442), .A1 (n_214), .B0 (latched_branch), .B1
       (n_6707), .Y (n_370));
  AOI22XL g180668(.A0 (n_442), .A1 (n_144), .B0 (latched_branch), .B1
       (n_6698), .Y (n_1514));
  AOI22XL g180669(.A0 (n_442), .A1 (n_146), .B0 (latched_branch), .B1
       (n_6699), .Y (n_1512));
  AO22X2 g180670(.A0 (n_442), .A1 (n_172), .B0 (latched_branch), .B1
       (n_6690), .Y (n_388));
  AO22X2 g180671(.A0 (n_442), .A1 (n_176), .B0 (latched_branch), .B1
       (n_6684), .Y (n_386));
  AO22X2 g180672(.A0 (n_442), .A1 (n_186), .B0 (latched_branch), .B1
       (n_6689), .Y (n_384));
  AO22X2 g180673(.A0 (n_442), .A1 (n_184), .B0 (latched_branch), .B1
       (n_6688), .Y (n_402));
  AO22X2 g180674(.A0 (n_442), .A1 (n_200), .B0 (latched_branch), .B1
       (n_6700), .Y (n_380));
  AO22X2 g180675(.A0 (n_442), .A1 (n_202), .B0 (latched_branch), .B1
       (n_6701), .Y (n_378));
  AO22X2 g180676(.A0 (n_442), .A1 (n_212), .B0 (latched_branch), .B1
       (n_6706), .Y (n_392));
  AO22X2 g180677(.A0 (n_442), .A1 (n_210), .B0 (latched_branch), .B1
       (n_6705), .Y (n_390));
  AO22X2 g180678(.A0 (n_442), .A1 (n_204), .B0 (latched_branch), .B1
       (n_6702), .Y (n_376));
  AO22X2 g180679(.A0 (n_442), .A1 (n_216), .B0 (latched_branch), .B1
       (n_6708), .Y (n_404));
  AO22X2 g180680(.A0 (n_442), .A1 (n_192), .B0 (latched_branch), .B1
       (n_6693), .Y (n_396));
  AO22X2 g180681(.A0 (n_442), .A1 (n_194), .B0 (latched_branch), .B1
       (n_6694), .Y (n_412));
  AO22X2 g180682(.A0 (n_442), .A1 (n_188), .B0 (latched_branch), .B1
       (n_6691), .Y (n_374));
  AO22X2 g180683(.A0 (n_442), .A1 (n_180), .B0 (latched_branch), .B1
       (n_6686), .Y (n_372));
  AO22X2 g180684(.A0 (n_442), .A1 (n_206), .B0 (latched_branch), .B1
       (n_6703), .Y (n_400));
  AO22X2 g180685(.A0 (n_442), .A1 (n_182), .B0 (latched_branch), .B1
       (n_6687), .Y (n_408));
  AO22X2 g180686(.A0 (n_442), .A1 (n_190), .B0 (latched_branch), .B1
       (n_6692), .Y (n_414));
  AO22X2 g180687(.A0 (n_442), .A1 (n_178), .B0 (latched_branch), .B1
       (n_6685), .Y (n_418));
  AO22X2 g180688(.A0 (n_442), .A1 (n_174), .B0 (latched_branch), .B1
       (n_6683), .Y (n_362));
  AO22X2 g180689(.A0 (n_442), .A1 (n_170), .B0 (latched_branch), .B1
       (n_6681), .Y (n_416));
  AO22X2 g180690(.A0 (n_442), .A1 (n_168), .B0 (latched_branch), .B1
       (n_6680), .Y (n_368));
  AO22X2 g180691(.A0 (n_442), .A1 (n_166), .B0 (latched_branch), .B1
       (n_6679), .Y (n_366));
  AO22X2 g180692(.A0 (n_442), .A1 (n_198), .B0 (latched_branch), .B1
       (n_6697), .Y (n_364));
  INVX1 g180693(.A (n_1369), .Y (n_1370));
  INVX1 g180694(.A (n_1366), .Y (n_1367));
  INVX1 g180696(.A (n_1343), .Y (n_1342));
  INVX1 g180700(.A (n_1330), .Y (n_1329));
  INVX1 g180701(.A (n_1328), .Y (n_1327));
  NAND2X1 g180708(.A (n_867), .B (n_858), .Y (n_1308));
  NAND2X1 g180709(.A (n_860), .B (n_861), .Y (n_1307));
  OAI21X1 g180710(.A0 (instr_lbu), .A1 (instr_lb), .B0 (cpu_state[0]),
       .Y (n_1306));
  OAI21X1 g180711(.A0 (\reg_op2[9]_9678 ), .A1 (\reg_op1[9]_9646 ), .B0
       (n_120), .Y (n_1305));
  NAND2X1 g180712(.A (decoded_rs2[1]), .B (n_953), .Y (n_1304));
  NAND2X1 g180713(.A (decoded_rs2[2]), .B (n_953), .Y (n_1303));
  OAI2BB1X1 g180714(.A0N (pcpi_timeout_counter[2]), .A1N (n_162), .B0
       (n_218), .Y (n_1302));
  OAI2BB1X1 g180715(.A0N (pcpi_timeout_counter[1]), .A1N
       (pcpi_timeout_counter[0]), .B0 (n_162), .Y (n_1301));
  AOI2BB1XL g180716(.A0N (latched_is_lu), .A1N (latched_is_lh), .B0
       (n_5984), .Y (n_1300));
  NAND2X1 g180717(.A (decoded_rs1[2]), .B (n_953), .Y (n_1299));
  NAND2X1 g180735(.A (decoded_rs1[0]), .B (n_953), .Y (n_1282));
  NAND2X1 g180736(.A (mem_rdata[5]), .B (n_839), .Y (n_1281));
  NAND2X1 g180737(.A (decoded_imm_j[14]), .B (n_953), .Y (n_1280));
  NAND2X1 g180739(.A (decoded_imm_j[18]), .B (n_953), .Y (n_1278));
  OAI21X1 g180745(.A0 (instr_lhu), .A1 (instr_lh), .B0 (cpu_state[0]),
       .Y (n_1272));
  NAND2X1 g180746(.A (mem_rdata[7]), .B (n_839), .Y (n_1271));
  NAND2X1 g180748(.A (decoded_imm_j[1]), .B (n_953), .Y (n_1269));
  OAI2BB1X1 g180750(.A0N (n_630), .A1N (n_628), .B0 (n_120), .Y
       (n_1267));
  NAND2X1 g180751(.A (decoded_imm_j[3]), .B (n_953), .Y (n_1266));
  NAND3X1 g180754(.A (\reg_op2[0]_9669 ), .B (reg_op1[0]), .C (n_283),
       .Y (n_1263));
  NAND2X1 g180756(.A (decoded_imm_j[4]), .B (n_953), .Y (n_1261));
  NAND2X1 g180758(.A (decoded_imm_j[2]), .B (n_953), .Y (n_1259));
  NAND2X1 g180759(.A (decoded_rd[2]), .B (n_953), .Y (n_1258));
  NAND2X1 g180761(.A (mem_rdata[6]), .B (n_839), .Y (n_1256));
  NAND2X1 g180763(.A (decoded_imm_j[20]), .B (n_953), .Y (n_1254));
  NAND3X1 g180769(.A (\reg_op1[20]_9657 ), .B
       (\genblk2.pcpi_div_minus_2470_59_n_500 ), .C (n_152), .Y
       (n_1248));
  NAND2X1 g180783(.A (mem_rdata[4]), .B (n_839), .Y (n_1234));
  NAND2X1 g180784(.A (decoded_imm_j[13]), .B (n_953), .Y (n_1233));
  NAND2X1 g180785(.A (decoded_rd[1]), .B (n_953), .Y (n_1232));
  NAND3BXL g180786(.AN (\genblk2.pcpi_div_quotient_msk [7]), .B
       (\genblk2.pcpi_div_running ), .C (n_734), .Y (n_1231));
  NOR2X1 g180804(.A (n_664), .B (n_150), .Y (n_1369));
  NOR2X1 g180805(.A (n_987), .B (n_573), .Y (n_1368));
  NOR2X1 g180806(.A (n_987), .B (n_627), .Y (n_1366));
  NOR2X1 g180808(.A (n_544), .B (n_668), .Y (n_1365));
  NOR2X1 g180809(.A (mem_rdata_latched[1]), .B (n_978), .Y (n_1364));
  NAND2X1 g180819(.A (n_991), .B (n_982), .Y (n_1363));
  AOI22X1 g180820(.A0 (mem_rdata_q[3]), .A1 (n_445), .B0
       (mem_rdata[3]), .B1 (n_446), .Y (n_1362));
  NAND3X1 g180822(.A (n_595), .B (n_833), .C (n_219), .Y (n_1361));
  NOR2BX1 g180823(.AN (n_870), .B (n_873), .Y (n_1360));
  NOR2BX1 g180838(.AN (n_863), .B (n_856), .Y (n_1359));
  NAND2X1 g180839(.A (n_857), .B (n_136), .Y (n_1358));
  NAND2X1 g180870(.A (n_652), .B (n_666), .Y (n_1357));
  NOR2X1 g180874(.A (cpu_state[6]), .B (n_849), .Y (n_1216));
  NOR3X1 g180875(.A (mem_rdata_q[23]), .B (mem_rdata_q[21]), .C
       (mem_rdata_q[22]), .Y (n_1356));
  NOR2X1 g180876(.A (cpu_state[2]), .B (n_833), .Y (n_1355));
  NAND2X1 g180877(.A (n_11740), .B (n_865), .Y (n_1354));
  NAND2X1 g180878(.A (n_3), .B (n_860), .Y (n_1353));
  NOR2BX1 g180879(.AN (n_855), .B (n_859), .Y (n_1352));
  NOR2BX1 g180881(.AN (n_984), .B (n_0), .Y (n_1351));
  AND2X1 g180883(.A (n_5), .B (n_3), .Y (n_1350));
  AND2X1 g180885(.A (n_871), .B (n_857), .Y (n_1349));
  NAND2X1 g180886(.A (n_11739), .B (n_869), .Y (n_1348));
  NAND2X1 g180887(.A (n_5), .B (n_861), .Y (n_1347));
  NAND2X1 g180888(.A (n_862), .B (n_867), .Y (n_1346));
  NAND2X1 g180890(.A (n_633), .B (n_988), .Y (n_1345));
  NOR2X1 g180891(.A (mem_rdata_q[12]), .B (n_877), .Y (n_1344));
  AND2X1 g180892(.A (n_977), .B (n_642), .Y (n_1343));
  OAI2BB1X1 g180893(.A0N (n_6532), .A1N (n_158), .B0 (n_545), .Y
       (n_1341));
  NOR2X1 g180894(.A (n_991), .B (n_854), .Y (n_1340));
  NOR3X1 g180896(.A (pcpi_div_wr), .B (pcpi_mul_wr), .C (pcpi_ready),
       .Y (n_1339));
  NOR2X1 g180897(.A (n_616), .B (n_877), .Y (n_1338));
  NOR2X1 g180898(.A (mem_rdata_q[12]), .B (n_874), .Y (n_1337));
  NAND2X1 g180899(.A (decoded_rs2[0]), .B (n_882), .Y (n_1336));
  NOR2X1 g180901(.A (decoded_rs2[0]), .B (n_880), .Y (n_1335));
  NAND2X1 g180904(.A (decoded_rs2[0]), .B (n_988), .Y (n_1334));
  NOR2X1 g180905(.A (decoded_rs2[0]), .B (n_885), .Y (n_1333));
  OR2X1 g180906(.A (n_633), .B (n_885), .Y (n_1332));
  NAND2X1 g180907(.A (n_587), .B (n_979), .Y (n_1331));
  NOR2X1 g180908(.A (n_974), .B (n_978), .Y (n_1330));
  NAND2X1 g180909(.A (n_851), .B (n_875), .Y (n_1328));
  NOR2X1 g180910(.A (mem_rdata_q[12]), .B (n_853), .Y (n_1326));
  NOR2X1 g180911(.A (n_616), .B (n_874), .Y (n_1325));
  NOR2BX1 g180913(.AN (n_976), .B (n_228), .Y (n_1324));
  AND2X1 g180914(.A (n_992), .B (n_616), .Y (n_1323));
  NOR3X1 g180915(.A (reg_sh[3]), .B (reg_sh[2]), .C (reg_sh[4]), .Y
       (n_1322));
  AND2X1 g180916(.A (n_992), .B (mem_rdata_q[12]), .Y (n_1321));
  NOR2BX1 g180917(.AN (n_976), .B (n_122), .Y (n_1320));
  OAI21X1 g180918(.A0 (n_613), .A1 (n_130), .B0 (n_324), .Y (n_1319));
  AND3XL g180919(.A (latched_is_lu), .B (cpu_state[0]), .C (n_608), .Y
       (n_1318));
  NAND2X2 g180920(.A (n_276), .B (n_667), .Y (n_335));
  OR2X1 g180921(.A (n_276), .B (n_953), .Y (n_342));
  AND2X1 g180922(.A (n_961), .B (cpu_state[5]), .Y (n_547));
  AND2X2 g180923(.A (decoder_trigger), .B (n_658), .Y (n_353));
  AND2X2 g180924(.A (n_820), .B (n_658), .Y (n_436));
  AND2X2 g180925(.A (n_980), .B (n_659), .Y (n_421));
  OR2X2 g180926(.A (n_664), .B (n_60), .Y (n_542));
  AND2X4 g180927(.A (n_773), .B (n_942), .Y (n_1310));
  AOI22XL g180928(.A0 (\genblk1.pcpi_mul_rd [34]), .A1 (n_11690), .B0
       (\genblk1.pcpi_mul_rd [2]), .B1 (n_59812_BAR), .Y (n_1192));
  NOR3BX1 g180929(.AN (n_320), .B (decoder_trigger), .C (n_324), .Y
       (n_1191));
  OAI2BB1X1 g180930(.A0N (n_14409_BAR), .A1N (n_96), .B0 (n_548), .Y
       (n_1190));
  OAI2BB1X1 g180932(.A0N (n_14409_BAR), .A1N (n_100), .B0 (n_548), .Y
       (n_1188));
  OAI2BB1X1 g180933(.A0N (n_14409_BAR), .A1N (n_110), .B0 (n_548), .Y
       (n_1187));
  OAI2BB1X1 g180934(.A0N (n_14409_BAR), .A1N (n_82), .B0 (n_548), .Y
       (n_1186));
  OAI2BB1X1 g180935(.A0N (n_14409_BAR), .A1N (n_104), .B0 (n_548), .Y
       (n_1185));
  OAI2BB1X1 g180936(.A0N (n_14409_BAR), .A1N (n_115), .B0 (n_548), .Y
       (n_1184));
  OAI2BB1X1 g180937(.A0N (n_14409_BAR), .A1N (n_84), .B0 (n_548), .Y
       (n_1183));
  OAI2BB1X1 g180938(.A0N (n_14409_BAR), .A1N (n_92), .B0 (n_548), .Y
       (n_1182));
  OAI2BB1X1 g180939(.A0N (n_14409_BAR), .A1N (n_94), .B0 (n_548), .Y
       (n_1181));
  OAI2BB1X1 g180942(.A0N (n_14409_BAR), .A1N (n_108), .B0 (n_548), .Y
       (n_1178));
  OAI2BB1X1 g180943(.A0N (n_14409_BAR), .A1N (n_90), .B0 (n_548), .Y
       (n_1177));
  OAI2BB1X1 g180944(.A0N (n_14409_BAR), .A1N (n_86), .B0 (n_548), .Y
       (n_1176));
  OAI2BB1X1 g180946(.A0N (n_14409_BAR), .A1N (n_98), .B0 (n_548), .Y
       (n_1174));
  OAI2BB1X1 g180947(.A0N (n_14409_BAR), .A1N (n_102), .B0 (n_548), .Y
       (n_1173));
  OAI2BB1X1 g180950(.A0N (n_14409_BAR), .A1N (n_88), .B0 (n_548), .Y
       (n_1170));
  OAI2BB1X1 g180951(.A0N (n_14409_BAR), .A1N (n_106), .B0 (n_548), .Y
       (n_1169));
  OAI2BB1X1 g180952(.A0N (n_14409_BAR), .A1N (n_112), .B0 (n_548), .Y
       (n_1168));
  MX2X1 g180953(.A (clear_prefetched_high_word_q), .B (n_222), .S0
       (n_6531), .Y (n_1167));
  AOI21X1 g180954(.A0 (last_mem_valid), .A1 (mem_la_firstword_reg), .B0
       (n_789), .Y (n_1166));
  OR4X1 g180955(.A (n_6672), .B (n_6674), .C (n_6660), .D (n_6658), .Y
       (n_1165));
  AOI22XL g180958(.A0 (pcpi_div_rd[20]), .A1 (n_39), .B0 (pcpi_rd[20]),
       .B1 (n_11689), .Y (n_1162));
  AOI22XL g180959(.A0 (pcpi_div_rd[21]), .A1 (n_39), .B0 (pcpi_rd[21]),
       .B1 (n_11689), .Y (n_1161));
  AOI22XL g180960(.A0 (pcpi_div_rd[22]), .A1 (n_39), .B0 (pcpi_rd[22]),
       .B1 (n_11689), .Y (n_1160));
  AOI22XL g180961(.A0 (pcpi_div_rd[31]), .A1 (n_39), .B0 (pcpi_rd[31]),
       .B1 (n_11689), .Y (n_1159));
  AOI22XL g180962(.A0 (pcpi_rd[2]), .A1 (n_11689), .B0
       (count_instr[34]), .B1 (instr_rdinstrh), .Y (n_1158));
  AOI22X1 g180963(.A0 (count_instr[56]), .A1 (instr_rdinstrh), .B0
       (count_instr[24]), .B1 (instr_rdinstr), .Y (n_1157));
  AOI22X1 g180964(.A0 (count_cycle[55]), .A1 (instr_rdcycleh), .B0
       (count_cycle[23]), .B1 (instr_rdcycle), .Y (n_1156));
  AOI22XL g180965(.A0 (\genblk1.pcpi_mul_rd [62]), .A1 (n_11690), .B0
       (\genblk1.pcpi_mul_rd [30]), .B1 (n_59812_BAR), .Y (n_1155));
  AOI22X1 g180966(.A0 (count_cycle[57]), .A1 (instr_rdcycleh), .B0
       (count_cycle[25]), .B1 (instr_rdcycle), .Y (n_1154));
  AOI22X1 g180967(.A0 (cpu_state[3]), .A1 (n_54), .B0 (count_instr[1]),
       .B1 (instr_rdinstr), .Y (n_1153));
  AOI22XL g180968(.A0 (\genblk1.pcpi_mul_rd [55]), .A1 (n_11690), .B0
       (\genblk1.pcpi_mul_rd [23]), .B1 (n_59812_BAR), .Y (n_1152));
  AOI22X1 g180969(.A0 (count_instr[55]), .A1 (instr_rdinstrh), .B0
       (count_instr[23]), .B1 (instr_rdinstr), .Y (n_1151));
  AOI22X1 g180970(.A0 (count_cycle[61]), .A1 (instr_rdcycleh), .B0
       (count_cycle[29]), .B1 (instr_rdcycle), .Y (n_1150));
  AOI22X1 g180971(.A0 (count_instr[53]), .A1 (instr_rdinstrh), .B0
       (count_instr[21]), .B1 (instr_rdinstr), .Y (n_1149));
  AOI22X1 g180972(.A0 (count_cycle[53]), .A1 (instr_rdcycleh), .B0
       (count_cycle[21]), .B1 (instr_rdcycle), .Y (n_1148));
  AOI22XL g180973(.A0 (pcpi_rd[17]), .A1 (n_11689), .B0
       (\genblk1.pcpi_mul_rd [17]), .B1 (n_59812_BAR), .Y (n_1147));
  AOI22X1 g180974(.A0 (count_instr[49]), .A1 (instr_rdinstrh), .B0
       (count_instr[17]), .B1 (instr_rdinstr), .Y (n_1146));
  AOI22X1 g180975(.A0 (count_instr[48]), .A1 (instr_rdinstrh), .B0
       (count_instr[16]), .B1 (instr_rdinstr), .Y (n_1145));
  AOI22XL g180976(.A0 (\genblk1.pcpi_mul_rd [60]), .A1 (n_11690), .B0
       (\genblk1.pcpi_mul_rd [28]), .B1 (n_59812_BAR), .Y (n_1144));
  AOI22X1 g180977(.A0 (count_cycle[48]), .A1 (instr_rdcycleh), .B0
       (count_cycle[16]), .B1 (instr_rdcycle), .Y (n_1143));
  AOI22XL g180978(.A0 (pcpi_div_rd[28]), .A1 (n_39), .B0 (pcpi_rd[28]),
       .B1 (n_11689), .Y (n_1142));
  AOI22X1 g180979(.A0 (count_instr[58]), .A1 (instr_rdinstrh), .B0
       (count_instr[26]), .B1 (instr_rdinstr), .Y (n_1141));
  AOI22X1 g180980(.A0 (count_cycle[60]), .A1 (instr_rdcycleh), .B0
       (count_cycle[28]), .B1 (instr_rdcycle), .Y (n_1140));
  AOI22XL g180981(.A0 (\genblk1.pcpi_mul_rd [38]), .A1 (n_11690), .B0
       (\genblk1.pcpi_mul_rd [6]), .B1 (n_59812_BAR), .Y (n_1139));
  AOI22X1 g180982(.A0 (count_cycle[47]), .A1 (instr_rdcycleh), .B0
       (count_cycle[15]), .B1 (instr_rdcycle), .Y (n_1138));
  AOI22XL g180983(.A0 (pcpi_div_rd[4]), .A1 (n_39), .B0
       (count_cycle[4]), .B1 (instr_rdcycle), .Y (n_1137));
  AOI22XL g180984(.A0 (pcpi_div_rd[26]), .A1 (n_39), .B0 (pcpi_rd[26]),
       .B1 (n_11689), .Y (n_1136));
  AOI22XL g180985(.A0 (pcpi_rd[4]), .A1 (n_11689), .B0
       (count_instr[36]), .B1 (instr_rdinstrh), .Y (n_1135));
  AOI22X1 g180986(.A0 (count_instr[54]), .A1 (instr_rdinstrh), .B0
       (count_instr[22]), .B1 (instr_rdinstr), .Y (n_1134));
  AOI22XL g180987(.A0 (\genblk1.pcpi_mul_rd [58]), .A1 (n_11690), .B0
       (\genblk1.pcpi_mul_rd [26]), .B1 (n_59812_BAR), .Y (n_1133));
  AOI22XL g180988(.A0 (\genblk1.pcpi_mul_rd [54]), .A1 (n_11690), .B0
       (\genblk1.pcpi_mul_rd [22]), .B1 (n_59812_BAR), .Y (n_1132));
  AOI22X1 g180989(.A0 (count_cycle[46]), .A1 (instr_rdcycleh), .B0
       (count_cycle[14]), .B1 (instr_rdcycle), .Y (n_1131));
  AOI22XL g180990(.A0 (pcpi_div_rd[14]), .A1 (n_39), .B0 (pcpi_rd[14]),
       .B1 (n_11689), .Y (n_1130));
  AOI22X1 g180991(.A0 (count_cycle[63]), .A1 (instr_rdcycleh), .B0
       (count_cycle[31]), .B1 (instr_rdcycle), .Y (n_1129));
  AOI22X1 g180992(.A0 (count_instr[46]), .A1 (instr_rdinstrh), .B0
       (count_instr[14]), .B1 (instr_rdinstr), .Y (n_1128));
  AOI22XL g180993(.A0 (pcpi_div_rd[9]), .A1 (n_39), .B0 (pcpi_rd[9]),
       .B1 (n_11689), .Y (n_1127));
  AOI22X1 g180994(.A0 (count_instr[51]), .A1 (instr_rdinstrh), .B0
       (count_instr[19]), .B1 (instr_rdinstr), .Y (n_1126));
  OAI22X1 g180995(.A0 (n_311), .A1 (n_601), .B0 (n_331), .B1 (n_653),
       .Y (n_1125));
  AOI22XL g180996(.A0 (\genblk1.pcpi_mul_rd [42]), .A1 (n_11690), .B0
       (\genblk1.pcpi_mul_rd [10]), .B1 (n_59812_BAR), .Y (n_1124));
  AOI22X1 g180997(.A0 (count_cycle[45]), .A1 (instr_rdcycleh), .B0
       (count_cycle[13]), .B1 (instr_rdcycle), .Y (n_1123));
  AOI22XL g180998(.A0 (\genblk1.pcpi_mul_rd [53]), .A1 (n_11690), .B0
       (\genblk1.pcpi_mul_rd [21]), .B1 (n_59812_BAR), .Y (n_1122));
  AOI22X1 g180999(.A0 (count_instr[45]), .A1 (instr_rdinstrh), .B0
       (count_instr[13]), .B1 (instr_rdinstr), .Y (n_1121));
  AOI22X1 g181000(.A0 (count_cycle[44]), .A1 (instr_rdcycleh), .B0
       (count_cycle[12]), .B1 (instr_rdcycle), .Y (n_1120));
  AOI22XL g181001(.A0 (pcpi_div_rd[18]), .A1 (n_39), .B0 (pcpi_rd[18]),
       .B1 (n_11689), .Y (n_1119));
  AOI22XL g181002(.A0 (pcpi_div_rd[12]), .A1 (n_39), .B0 (pcpi_rd[12]),
       .B1 (n_11689), .Y (n_1118));
  AOI22X1 g181003(.A0 (count_instr[44]), .A1 (instr_rdinstrh), .B0
       (count_instr[12]), .B1 (instr_rdinstr), .Y (n_1117));
  AOI22X1 g181004(.A0 (count_cycle[50]), .A1 (instr_rdcycleh), .B0
       (count_cycle[18]), .B1 (instr_rdcycle), .Y (n_1116));
  AOI22X1 g181005(.A0 (count_instr[52]), .A1 (instr_rdinstrh), .B0
       (count_instr[20]), .B1 (instr_rdinstr), .Y (n_1115));
  AOI22X1 g181006(.A0 (count_instr[59]), .A1 (instr_rdinstrh), .B0
       (count_instr[27]), .B1 (instr_rdinstr), .Y (n_1114));
  AOI22XL g181007(.A0 (\genblk1.pcpi_mul_rd [44]), .A1 (n_11690), .B0
       (\genblk1.pcpi_mul_rd [12]), .B1 (n_59812_BAR), .Y (n_1113));
  AOI22X1 g181008(.A0 (count_cycle[41]), .A1 (instr_rdcycleh), .B0
       (count_cycle[9]), .B1 (instr_rdcycle), .Y (n_1112));
  AOI22XL g181009(.A0 (pcpi_div_rd[29]), .A1 (n_39), .B0 (pcpi_rd[29]),
       .B1 (n_11689), .Y (n_1111));
  AOI22X1 g181010(.A0 (count_cycle[56]), .A1 (instr_rdcycleh), .B0
       (count_cycle[24]), .B1 (instr_rdcycle), .Y (n_1110));
  AOI22XL g181011(.A0 (\genblk1.pcpi_mul_rd [50]), .A1 (n_11690), .B0
       (\genblk1.pcpi_mul_rd [18]), .B1 (n_59812_BAR), .Y (n_1109));
  AOI22XL g181012(.A0 (pcpi_div_rd[17]), .A1 (n_39), .B0
       (\genblk1.pcpi_mul_rd [49]), .B1 (n_11690), .Y (n_1108));
  AOI22X1 g181013(.A0 (count_cycle[58]), .A1 (instr_rdcycleh), .B0
       (count_cycle[26]), .B1 (instr_rdcycle), .Y (n_1107));
  AOI22XL g181014(.A0 (pcpi_div_rd[15]), .A1 (n_39), .B0 (pcpi_rd[15]),
       .B1 (n_11689), .Y (n_1106));
  AOI22XL g181015(.A0 (\genblk1.pcpi_mul_rd [46]), .A1 (n_11690), .B0
       (\genblk1.pcpi_mul_rd [14]), .B1 (n_59812_BAR), .Y (n_1105));
  AOI22XL g181016(.A0 (pcpi_div_rd[13]), .A1 (n_39), .B0 (pcpi_rd[13]),
       .B1 (n_11689), .Y (n_1104));
  AOI22XL g181017(.A0 (\genblk1.pcpi_mul_rd [45]), .A1 (n_11690), .B0
       (\genblk1.pcpi_mul_rd [13]), .B1 (n_59812_BAR), .Y (n_1103));
  AOI22XL g181018(.A0 (\genblk1.pcpi_mul_rd [3]), .A1 (n_59812_BAR),
       .B0 (count_cycle[3]), .B1 (instr_rdcycle), .Y (n_1102));
  AOI22X1 g181019(.A0 (count_instr[42]), .A1 (instr_rdinstrh), .B0
       (count_instr[10]), .B1 (instr_rdinstr), .Y (n_1101));
  AOI22XL g181020(.A0 (pcpi_div_rd[1]), .A1 (n_39), .B0 (pcpi_rd[1]),
       .B1 (n_11689), .Y (n_1100));
  AOI22X1 g181021(.A0 (count_instr[41]), .A1 (instr_rdinstrh), .B0
       (count_instr[9]), .B1 (instr_rdinstr), .Y (n_1099));
  AOI22X1 g181022(.A0 (count_instr[47]), .A1 (instr_rdinstrh), .B0
       (count_instr[15]), .B1 (instr_rdinstr), .Y (n_1098));
  AOI22XL g181023(.A0 (\genblk1.pcpi_mul_rd [61]), .A1 (n_11690), .B0
       (\genblk1.pcpi_mul_rd [29]), .B1 (n_59812_BAR), .Y (n_1097));
  AOI22X1 g181024(.A0 (count_instr[39]), .A1 (instr_rdinstrh), .B0
       (count_instr[7]), .B1 (instr_rdinstr), .Y (n_1096));
  AOI22XL g181025(.A0 (\genblk1.pcpi_mul_rd [39]), .A1 (n_11690), .B0
       (\genblk1.pcpi_mul_rd [7]), .B1 (n_59812_BAR), .Y (n_1095));
  OAI22X1 g181026(.A0 (n_343), .A1 (n_656), .B0 (n_331), .B1 (n_598),
       .Y (n_1094));
  AOI22XL g181027(.A0 (pcpi_div_rd[6]), .A1 (n_39), .B0 (pcpi_rd[6]),
       .B1 (n_11689), .Y (n_1093));
  AOI22X1 g181028(.A0 (count_cycle[38]), .A1 (instr_rdcycleh), .B0
       (count_cycle[6]), .B1 (instr_rdcycle), .Y (n_1092));
  AOI22XL g181029(.A0 (\genblk1.pcpi_mul_rd [48]), .A1 (n_11690), .B0
       (\genblk1.pcpi_mul_rd [16]), .B1 (n_59812_BAR), .Y (n_1091));
  AOI22XL g181030(.A0 (pcpi_div_rd[5]), .A1 (n_39), .B0 (pcpi_rd[5]),
       .B1 (n_11689), .Y (n_1090));
  AOI22X1 g181031(.A0 (count_instr[38]), .A1 (instr_rdinstrh), .B0
       (count_instr[6]), .B1 (instr_rdinstr), .Y (n_1089));
  AOI22XL g181032(.A0 (\genblk1.pcpi_mul_rd [37]), .A1 (n_11690), .B0
       (\genblk1.pcpi_mul_rd [5]), .B1 (n_59812_BAR), .Y (n_1088));
  AOI22X1 g181033(.A0 (count_instr[4]), .A1 (instr_rdinstr), .B0
       (count_cycle[36]), .B1 (instr_rdcycleh), .Y (n_1087));
  AOI22X1 g181034(.A0 (count_instr[40]), .A1 (instr_rdinstrh), .B0
       (count_instr[8]), .B1 (instr_rdinstr), .Y (n_1086));
  AOI22X1 g181035(.A0 (count_instr[61]), .A1 (instr_rdinstrh), .B0
       (count_instr[29]), .B1 (instr_rdinstr), .Y (n_1085));
  AOI22XL g181036(.A0 (pcpi_rd[3]), .A1 (n_11689), .B0
       (\genblk1.pcpi_mul_rd [35]), .B1 (n_11690), .Y (n_1084));
  AOI22X1 g181037(.A0 (count_instr[3]), .A1 (instr_rdinstr), .B0
       (count_cycle[35]), .B1 (instr_rdcycleh), .Y (n_1083));
  AOI22X1 g181038(.A0 (count_cycle[59]), .A1 (instr_rdcycleh), .B0
       (count_cycle[27]), .B1 (instr_rdcycle), .Y (n_1082));
  AOI22X1 g181039(.A0 (mem_rdata_q[15]), .A1 (n_712), .B0
       (mem_rdata[15]), .B1 (n_745), .Y (n_1081));
  AOI22X1 g181040(.A0 (count_instr[2]), .A1 (instr_rdinstr), .B0
       (count_cycle[34]), .B1 (instr_rdcycleh), .Y (n_1080));
  AOI22X1 g181041(.A0 (count_instr[37]), .A1 (instr_rdinstrh), .B0
       (count_instr[5]), .B1 (instr_rdinstr), .Y (n_1079));
  AOI22X1 g181042(.A0 (count_cycle[43]), .A1 (instr_rdcycleh), .B0
       (count_cycle[11]), .B1 (instr_rdcycle), .Y (n_1078));
  AOI22X1 g181043(.A0 (count_instr[57]), .A1 (instr_rdinstrh), .B0
       (count_instr[25]), .B1 (instr_rdinstr), .Y (n_1077));
  AOI22XL g181044(.A0 (\genblk1.pcpi_mul_rd [1]), .A1 (n_59812_BAR),
       .B0 (count_instr[33]), .B1 (instr_rdinstrh), .Y (n_1076));
  AOI22XL g181045(.A0 (pcpi_div_rd[2]), .A1 (n_39), .B0
       (count_cycle[2]), .B1 (instr_rdcycle), .Y (n_1075));
  AOI22X1 g181046(.A0 (count_cycle[37]), .A1 (instr_rdcycleh), .B0
       (count_cycle[5]), .B1 (instr_rdcycle), .Y (n_1074));
  AOI22XL g181047(.A0 (pcpi_rd[11]), .A1 (n_11689), .B0
       (\genblk1.pcpi_mul_rd [11]), .B1 (n_59812_BAR), .Y (n_1073));
  AOI22XL g181048(.A0 (pcpi_div_rd[3]), .A1 (n_39), .B0
       (count_instr[35]), .B1 (instr_rdinstrh), .Y (n_1072));
  AOI22X1 g181049(.A0 (count_cycle[49]), .A1 (instr_rdcycleh), .B0
       (count_cycle[17]), .B1 (instr_rdcycle), .Y (n_1071));
  AOI22XL g181050(.A0 (\genblk1.pcpi_mul_rd [59]), .A1 (n_11690), .B0
       (\genblk1.pcpi_mul_rd [27]), .B1 (n_59812_BAR), .Y (n_1070));
  AOI22X1 g181051(.A0 (count_cycle[40]), .A1 (instr_rdcycleh), .B0
       (count_cycle[8]), .B1 (instr_rdcycle), .Y (n_1069));
  AOI22X1 g181052(.A0 (count_instr[63]), .A1 (instr_rdinstrh), .B0
       (count_instr[31]), .B1 (instr_rdinstr), .Y (n_1068));
  AOI22XL g181053(.A0 (\genblk1.pcpi_mul_rd [41]), .A1 (n_11690), .B0
       (\genblk1.pcpi_mul_rd [9]), .B1 (n_59812_BAR), .Y (n_1067));
  AOI22X1 g181054(.A0 (count_instr[62]), .A1 (instr_rdinstrh), .B0
       (count_instr[30]), .B1 (instr_rdinstr), .Y (n_1066));
  AOI22X1 g181055(.A0 (count_cycle[39]), .A1 (instr_rdcycleh), .B0
       (count_cycle[7]), .B1 (instr_rdcycle), .Y (n_1065));
  AOI22X1 g181056(.A0 (count_cycle[42]), .A1 (instr_rdcycleh), .B0
       (count_cycle[10]), .B1 (instr_rdcycle), .Y (n_1064));
  AOI22X1 g181057(.A0 (count_cycle[62]), .A1 (instr_rdcycleh), .B0
       (count_cycle[30]), .B1 (instr_rdcycle), .Y (n_1063));
  AOI22XL g181058(.A0 (pcpi_div_rd[16]), .A1 (n_39), .B0 (pcpi_rd[16]),
       .B1 (n_11689), .Y (n_1062));
  AOI22XL g181059(.A0 (pcpi_div_rd[27]), .A1 (n_39), .B0 (pcpi_rd[27]),
       .B1 (n_11689), .Y (n_1061));
  AOI22X1 g181060(.A0 (count_cycle[54]), .A1 (instr_rdcycleh), .B0
       (count_cycle[22]), .B1 (instr_rdcycle), .Y (n_1060));
  AOI22XL g181061(.A0 (\genblk1.pcpi_mul_rd [56]), .A1 (n_11690), .B0
       (\genblk1.pcpi_mul_rd [24]), .B1 (n_59812_BAR), .Y (n_1059));
  AOI22XL g181062(.A0 (\genblk1.pcpi_mul_rd [36]), .A1 (n_11690), .B0
       (\genblk1.pcpi_mul_rd [4]), .B1 (n_59812_BAR), .Y (n_1058));
  AOI22XL g181063(.A0 (pcpi_div_rd[7]), .A1 (n_39), .B0 (pcpi_rd[7]),
       .B1 (n_11689), .Y (n_1057));
  AOI22XL g181064(.A0 (\genblk1.pcpi_mul_rd [47]), .A1 (n_11690), .B0
       (\genblk1.pcpi_mul_rd [15]), .B1 (n_59812_BAR), .Y (n_1056));
  AOI22X1 g181065(.A0 (count_cycle[52]), .A1 (instr_rdcycleh), .B0
       (count_cycle[20]), .B1 (instr_rdcycle), .Y (n_1055));
  AOI22XL g181066(.A0 (pcpi_div_rd[24]), .A1 (n_39), .B0 (pcpi_rd[24]),
       .B1 (n_11689), .Y (n_1054));
  AOI22XL g181067(.A0 (\genblk1.pcpi_mul_rd [51]), .A1 (n_11690), .B0
       (\genblk1.pcpi_mul_rd [19]), .B1 (n_59812_BAR), .Y (n_1053));
  AOI22X1 g181068(.A0 (count_instr[60]), .A1 (instr_rdinstrh), .B0
       (count_instr[28]), .B1 (instr_rdinstr), .Y (n_1052));
  AOI22XL g181069(.A0 (\genblk1.pcpi_mul_rd [52]), .A1 (n_11690), .B0
       (\genblk1.pcpi_mul_rd [20]), .B1 (n_59812_BAR), .Y (n_1051));
  AOI22XL g181070(.A0 (\genblk1.pcpi_mul_rd [57]), .A1 (n_11690), .B0
       (\genblk1.pcpi_mul_rd [25]), .B1 (n_59812_BAR), .Y (n_1050));
  AOI22XL g181071(.A0 (pcpi_div_rd[30]), .A1 (n_39), .B0 (pcpi_rd[30]),
       .B1 (n_11689), .Y (n_1049));
  AOI22XL g181072(.A0 (\genblk1.pcpi_mul_rd [63]), .A1 (n_11690), .B0
       (\genblk1.pcpi_mul_rd [31]), .B1 (n_59812_BAR), .Y (n_1048));
  AOI22XL g181073(.A0 (pcpi_div_rd[8]), .A1 (n_39), .B0 (pcpi_rd[8]),
       .B1 (n_11689), .Y (n_1047));
  AOI22XL g181074(.A0 (pcpi_div_rd[10]), .A1 (n_39), .B0 (pcpi_rd[10]),
       .B1 (n_11689), .Y (n_1046));
  AOI22X1 g181075(.A0 (count_instr[43]), .A1 (instr_rdinstrh), .B0
       (count_instr[11]), .B1 (instr_rdinstr), .Y (n_1045));
  AOI22XL g181076(.A0 (pcpi_div_rd[11]), .A1 (n_39), .B0
       (\genblk1.pcpi_mul_rd [43]), .B1 (n_11690), .Y (n_1044));
  AOI22XL g181077(.A0 (\genblk1.pcpi_mul_rd [40]), .A1 (n_11690), .B0
       (\genblk1.pcpi_mul_rd [8]), .B1 (n_59812_BAR), .Y (n_1043));
  AOI22XL g181078(.A0 (pcpi_div_rd[23]), .A1 (n_39), .B0 (pcpi_rd[23]),
       .B1 (n_11689), .Y (n_1042));
  AOI22X1 g181079(.A0 (count_instr[50]), .A1 (instr_rdinstrh), .B0
       (count_instr[18]), .B1 (instr_rdinstr), .Y (n_1041));
  AOI22X1 g181080(.A0 (count_cycle[51]), .A1 (instr_rdcycleh), .B0
       (count_cycle[19]), .B1 (instr_rdcycle), .Y (n_1040));
  AOI22XL g181081(.A0 (pcpi_div_rd[19]), .A1 (n_39), .B0 (pcpi_rd[19]),
       .B1 (n_11689), .Y (n_1039));
  AOI22XL g181082(.A0 (pcpi_div_rd[25]), .A1 (n_39), .B0 (pcpi_rd[25]),
       .B1 (n_11689), .Y (n_1038));
  AOI22X1 g181083(.A0 (mem_rdata_q[2]), .A1 (n_712), .B0
       (mem_rdata[2]), .B1 (n_745), .Y (n_1037));
  AOI22X1 g181084(.A0 (mem_rdata_q[5]), .A1 (n_712), .B0
       (mem_rdata[5]), .B1 (n_745), .Y (n_1036));
  AOI22X1 g181085(.A0 (mem_rdata_q[8]), .A1 (n_712), .B0
       (mem_rdata[8]), .B1 (n_745), .Y (n_1035));
  AOI22X1 g181086(.A0 (mem_rdata_q[9]), .A1 (n_712), .B0
       (mem_rdata[9]), .B1 (n_745), .Y (n_1034));
  AOI22X1 g181087(.A0 (mem_rdata_q[10]), .A1 (n_712), .B0
       (mem_rdata[10]), .B1 (n_745), .Y (n_1033));
  AOI22X1 g181088(.A0 (mem_rdata_q[11]), .A1 (n_712), .B0
       (mem_rdata[11]), .B1 (n_745), .Y (n_1032));
  AOI22X1 g181089(.A0 (mem_rdata_q[6]), .A1 (n_712), .B0
       (mem_rdata[6]), .B1 (n_745), .Y (n_1031));
  AOI22X1 g181090(.A0 (mem_rdata_q[4]), .A1 (n_712), .B0
       (mem_rdata[4]), .B1 (n_745), .Y (n_1030));
  AOI22X1 g181091(.A0 (mem_rdata_q[7]), .A1 (n_712), .B0
       (mem_rdata[7]), .B1 (n_745), .Y (n_1029));
  AOI22X1 g181092(.A0 (mem_rdata_q[12]), .A1 (n_712), .B0
       (mem_rdata[12]), .B1 (n_745), .Y (n_1028));
  MX2X1 g181093(.A (mem_rdata_q[1]), .B (mem_rdata_latched[1]), .S0
       (n_446), .Y (n_1027));
  MX2X1 g181094(.A (n_5613), .B (mem_rdata_q[28]), .S0 (n_538), .Y
       (n_1026));
  MX2X1 g181095(.A (n_5597), .B (mem_rdata_q[12]), .S0 (n_538), .Y
       (n_1025));
  MX2X1 g181096(.A (n_5595), .B (mem_rdata_q[10]), .S0 (n_538), .Y
       (n_1024));
  MX2X1 g181097(.A (n_5593), .B (mem_rdata_q[8]), .S0 (n_538), .Y
       (n_1023));
  MX2X1 g181098(.A (n_5585), .B (mem_rdata_q[0]), .S0 (n_538), .Y
       (n_1022));
  MX2X1 g181099(.A (n_5586), .B (mem_rdata_q[1]), .S0 (n_538), .Y
       (n_1021));
  MX2X1 g181100(.A (n_5588), .B (mem_rdata_q[3]), .S0 (n_538), .Y
       (n_1020));
  MX2X1 g181101(.A (n_5590), .B (mem_rdata_q[5]), .S0 (n_538), .Y
       (n_1019));
  MX2X1 g181102(.A (n_5591), .B (mem_rdata_q[6]), .S0 (n_538), .Y
       (n_1018));
  MX2X1 g181103(.A (n_5592), .B (mem_rdata_q[7]), .S0 (n_538), .Y
       (n_1017));
  MX2X1 g181104(.A (n_5594), .B (mem_rdata_q[9]), .S0 (n_538), .Y
       (n_1016));
  MX2X1 g181105(.A (n_5596), .B (mem_rdata_q[11]), .S0 (n_538), .Y
       (n_1015));
  MX2X1 g181106(.A (n_5598), .B (mem_rdata_q[13]), .S0 (n_538), .Y
       (n_1014));
  MX2X1 g181107(.A (n_5599), .B (mem_rdata_q[14]), .S0 (n_538), .Y
       (n_1013));
  MX2X1 g181108(.A (n_5600), .B (mem_rdata_q[15]), .S0 (n_538), .Y
       (n_1012));
  MX2X1 g181109(.A (n_5602), .B (mem_rdata_q[17]), .S0 (n_538), .Y
       (n_1011));
  MX2X1 g181110(.A (n_5603), .B (mem_rdata_q[18]), .S0 (n_538), .Y
       (n_1010));
  MX2X1 g181111(.A (n_5604), .B (mem_rdata_q[19]), .S0 (n_538), .Y
       (n_1009));
  MX2X1 g181112(.A (n_5606), .B (mem_rdata_q[21]), .S0 (n_538), .Y
       (n_1008));
  MX2X1 g181113(.A (n_5607), .B (mem_rdata_q[22]), .S0 (n_538), .Y
       (n_1007));
  MX2X1 g181114(.A (n_5608), .B (mem_rdata_q[23]), .S0 (n_538), .Y
       (n_1006));
  MX2X1 g181115(.A (n_5610), .B (mem_rdata_q[25]), .S0 (n_538), .Y
       (n_1005));
  MX2X1 g181116(.A (n_5612), .B (mem_rdata_q[27]), .S0 (n_538), .Y
       (n_1004));
  MX2X1 g181117(.A (n_5614), .B (mem_rdata_q[29]), .S0 (n_538), .Y
       (n_1003));
  MX2X1 g181118(.A (n_5615), .B (mem_rdata_q[30]), .S0 (n_538), .Y
       (n_1002));
  MX2X1 g181119(.A (n_5616), .B (mem_rdata_q[31]), .S0 (n_538), .Y
       (n_1001));
  MX2X1 g181120(.A (n_5605), .B (mem_rdata_q[20]), .S0 (n_538), .Y
       (n_1000));
  MX2X1 g181121(.A (n_5589), .B (mem_rdata_q[4]), .S0 (n_538), .Y
       (n_999));
  MX2X1 g181122(.A (n_5587), .B (mem_rdata_q[2]), .S0 (n_538), .Y
       (n_998));
  MX2X1 g181123(.A (n_5611), .B (mem_rdata_q[26]), .S0 (n_538), .Y
       (n_997));
  MX2X1 g181124(.A (n_5609), .B (mem_rdata_q[24]), .S0 (n_538), .Y
       (n_996));
  MX2X1 g181125(.A (n_5601), .B (mem_rdata_q[16]), .S0 (n_538), .Y
       (n_995));
  OAI22X1 g181126(.A0 (n_759), .A1 (n_446), .B0 (n_445), .B1 (n_345),
       .Y (n_994));
  NAND3BXL g181127(.AN (mem_rdata_q[3]), .B (mem_rdata_q[1]), .C
       (n_763), .Y (n_1215));
  AOI22X1 g181128(.A0 (mem_rdata_q[19]), .A1 (n_445), .B0
       (mem_rdata[19]), .B1 (n_446), .Y (n_1214));
  AOI22X1 g181129(.A0 (mem_rdata_q[23]), .A1 (n_445), .B0
       (mem_rdata[23]), .B1 (n_446), .Y (n_1213));
  AOI22X1 g181130(.A0 (mem_rdata_q[24]), .A1 (n_445), .B0
       (mem_rdata[24]), .B1 (n_446), .Y (n_1212));
  AOI22X1 g181131(.A0 (mem_rdata_q[21]), .A1 (n_445), .B0
       (mem_rdata[21]), .B1 (n_446), .Y (n_1211));
  AOI22X1 g181132(.A0 (mem_rdata_q[25]), .A1 (n_445), .B0
       (mem_rdata[25]), .B1 (n_446), .Y (n_1210));
  AOI22X1 g181133(.A0 (mem_rdata_q[18]), .A1 (n_445), .B0
       (mem_rdata[18]), .B1 (n_446), .Y (n_1209));
  AOI22X1 g181134(.A0 (mem_rdata_q[30]), .A1 (n_445), .B0
       (mem_rdata[30]), .B1 (n_446), .Y (n_1208));
  MX2X1 g181135(.A (mem_rdata[28]), .B (mem_rdata_q[28]), .S0 (n_445),
       .Y (n_1207));
  AOI22X1 g181136(.A0 (mem_rdata_q[22]), .A1 (n_445), .B0
       (mem_rdata[22]), .B1 (n_446), .Y (n_1206));
  MX2X1 g181137(.A (mem_rdata[27]), .B (mem_rdata_q[27]), .S0 (n_445),
       .Y (n_1205));
  AOI22X1 g181138(.A0 (mem_rdata_q[13]), .A1 (n_445), .B0
       (mem_rdata[13]), .B1 (n_446), .Y (n_1204));
  MX2X1 g181139(.A (mem_rdata[26]), .B (mem_rdata_q[26]), .S0 (n_445),
       .Y (n_1203));
  AOI22X1 g181140(.A0 (mem_rdata_q[20]), .A1 (n_445), .B0
       (mem_rdata[20]), .B1 (n_446), .Y (n_1202));
  AOI22X1 g181141(.A0 (mem_rdata_q[29]), .A1 (n_445), .B0
       (mem_rdata[29]), .B1 (n_446), .Y (n_1201));
  AOI22X1 g181142(.A0 (mem_rdata_q[31]), .A1 (n_445), .B0
       (mem_rdata[31]), .B1 (n_446), .Y (n_1200));
  OAI22X1 g181143(.A0 (n_228), .A1 (n_598), .B0 (n_122), .B1 (n_600),
       .Y (n_1199));
  OAI22X1 g181144(.A0 (\reg_op2[1]_9670 ), .A1 (n_565), .B0
       (\reg_op1[1]_9638 ), .B1 (n_629), .Y (n_1198));
  AOI22X1 g181145(.A0 (mem_rdata_q[14]), .A1 (n_445), .B0
       (mem_rdata[14]), .B1 (n_446), .Y (n_1197));
  AOI21X1 g181146(.A0 (\reg_op1[8]_9645 ), .A1
       (\genblk2.pcpi_div_minus_2470_59_n_492 ), .B0 (n_883), .Y
       (n_1196));
  AOI21X1 g181147(.A0 (\reg_op1[9]_9646 ), .A1 (n_714), .B0 (n_879), .Y
       (n_1195));
  AOI21X1 g181148(.A0 (reg_op1[0]), .A1 (n_630), .B0 (n_878), .Y
       (n_1194));
  NAND3X1 g181149(.A (mem_state[0]), .B (n_603), .C (n_446), .Y
       (n_1193));
  INVX1 g181150(.A (n_981), .Y (n_980));
  INVX1 g181151(.A (n_968), .Y (n_969));
  INVX1 g181152(.A (n_966), .Y (n_965));
  INVX1 g181153(.A (n_963), .Y (n_962));
  AND2X1 g181160(.A (n_6756), .B (n_543), .Y (n_951));
  AND2X1 g181161(.A (n_6749), .B (n_543), .Y (n_950));
  NAND2X1 g181162(.A (decoded_imm[24]), .B (n_537), .Y (n_949));
  AND2X1 g181163(.A (n_543), .B (n_6744), .Y (n_948));
  NOR2X1 g181164(.A (\reg_op2[1]_9670 ), .B (\reg_op1[1]_9638 ), .Y
       (n_947));
  AND2X1 g181165(.A (n_543), .B (n_6741), .Y (n_946));
  NAND2X1 g181166(.A (decoded_imm[22]), .B (n_537), .Y (n_945));
  AND2X1 g181167(.A (n_6784), .B (n_543), .Y (n_944));
  AND2X1 g181168(.A (n_6761), .B (n_543), .Y (n_943));
  NOR2XL g181169(.A (\genblk1.pcpi_mul_active [0]), .B (n_6565), .Y
       (n_942));
  AND2X1 g181170(.A (n_6794), .B (n_543), .Y (n_941));
  NOR2X1 g181171(.A (\reg_op2[14]_9683 ), .B (\reg_op1[14]_9651 ), .Y
       (n_940));
  AND2X1 g181172(.A (n_6752), .B (n_543), .Y (n_939));
  AND2X1 g181173(.A (n_6763), .B (n_543), .Y (n_938));
  NOR2X1 g181174(.A (\reg_op2[15]_9684 ), .B (\reg_op1[15]_9652 ), .Y
       (n_937));
  NAND2X1 g181175(.A (decoded_imm[25]), .B (n_537), .Y (n_936));
  NAND2X1 g181176(.A (mem_16bit_buffer[8]), .B (n_360), .Y (n_935));
  AND2X1 g181177(.A (n_6780), .B (n_543), .Y (n_934));
  AND2X1 g181178(.A (n_6774), .B (n_543), .Y (n_933));
  AND2X1 g181179(.A (n_6786), .B (n_543), .Y (n_932));
  NOR2BX1 g181180(.AN (latched_is_lu), .B (n_56), .Y (n_931));
  NAND2X1 g181181(.A (mem_16bit_buffer[5]), .B (n_360), .Y (n_930));
  AND2X1 g181182(.A (n_6793), .B (n_543), .Y (n_929));
  AND2X1 g181183(.A (n_6800), .B (n_543), .Y (n_928));
  AND2X1 g181184(.A (n_6764), .B (n_543), .Y (n_927));
  AND2X1 g181185(.A (n_6799), .B (n_543), .Y (n_926));
  AND2X1 g181186(.A (n_543), .B (n_6743), .Y (n_925));
  AND2X1 g181187(.A (n_6751), .B (n_543), .Y (n_924));
  NAND2X1 g181188(.A (decoded_imm[31]), .B (n_537), .Y (n_923));
  AND2X1 g181189(.A (n_6773), .B (n_543), .Y (n_922));
  NAND2X1 g181190(.A (mem_16bit_buffer[3]), .B (n_360), .Y (n_921));
  AND2X1 g181191(.A (n_6777), .B (n_543), .Y (n_920));
  AND2X1 g181192(.A (n_6778), .B (n_543), .Y (n_919));
  AND2X1 g181193(.A (n_6765), .B (n_543), .Y (n_918));
  NAND2XL g181194(.A (pcpi_wr), .B (n_11689), .Y (n_917));
  NOR2X1 g181195(.A (\reg_op2[8]_9677 ), .B (\reg_op1[8]_9645 ), .Y
       (n_916));
  NAND2X1 g181196(.A (mem_16bit_buffer[14]), .B (n_360), .Y (n_915));
  NOR2X1 g181197(.A (\reg_op2[6]_9675 ), .B (\reg_op1[6]_9643 ), .Y
       (n_914));
  AND2X1 g181198(.A (n_6791), .B (n_543), .Y (n_913));
  AND2X1 g181199(.A (n_6789), .B (n_543), .Y (n_912));
  NAND2X1 g181200(.A (decoded_imm[30]), .B (n_537), .Y (n_911));
  AND2X1 g181201(.A (n_6758), .B (n_543), .Y (n_910));
  AND2X1 g181202(.A (n_6790), .B (n_543), .Y (n_909));
  AND2X1 g181203(.A (n_6779), .B (n_543), .Y (n_908));
  AND2X1 g181204(.A (n_6802), .B (n_543), .Y (n_907));
  NAND2X1 g181205(.A (decoded_imm[28]), .B (n_537), .Y (n_906));
  NOR2X1 g181206(.A (mem_state[0]), .B (n_603), .Y (n_905));
  AND2X1 g181207(.A (n_6775), .B (n_543), .Y (n_904));
  NAND2X1 g181208(.A (decoded_imm[20]), .B (n_537), .Y (n_903));
  AND2X1 g181209(.A (n_6759), .B (n_543), .Y (n_902));
  NAND2X1 g181210(.A (prefetched_high_word), .B
       (clear_prefetched_high_word_q), .Y (n_901));
  NOR2X1 g181211(.A (\reg_op2[12]_9681 ), .B (\reg_op1[12]_9649 ), .Y
       (n_900));
  AND2X1 g181212(.A (n_6771), .B (n_543), .Y (n_899));
  AND2X1 g181213(.A (n_6753), .B (n_543), .Y (n_898));
  NOR2X1 g181214(.A (\reg_op2[7]_9676 ), .B (\reg_op1[7]_9644 ), .Y
       (n_897));
  NOR2X1 g181215(.A (count_cycle[0]), .B (n_544), .Y (n_896));
  AND2X1 g181216(.A (n_6768), .B (n_543), .Y (n_895));
  AND2X1 g181217(.A (n_6750), .B (n_543), .Y (n_894));
  AND2X1 g181218(.A (n_6770), .B (n_543), .Y (n_893));
  NAND2X1 g181219(.A (mem_16bit_buffer[13]), .B (n_360), .Y (n_892));
  AND2X1 g181220(.A (n_6801), .B (n_543), .Y (n_891));
  AND2X1 g181221(.A (n_543), .B (cpu_state[7]), .Y (n_890));
  AND2X1 g181222(.A (n_6767), .B (n_543), .Y (n_889));
  AND2X1 g181223(.A (n_6754), .B (n_543), .Y (n_888));
  NAND2X1 g181224(.A (decoded_imm[23]), .B (n_537), .Y (n_887));
  AND2X1 g181225(.A (n_6788), .B (n_543), .Y (n_886));
  OR2X1 g181226(.A (instr_slli), .B (instr_sll), .Y (n_993));
  NOR2X1 g181227(.A (mem_rdata_q[14]), .B (mem_rdata_q[13]), .Y
       (n_992));
  NOR2X1 g181228(.A (instr_srai), .B (instr_sra), .Y (n_991));
  NOR2BX1 g181229(.AN (latched_is_lh), .B (n_122), .Y (n_990));
  NAND2X1 g181230(.A (n_5617), .B (n_543), .Y (n_989));
  NOR2X1 g181231(.A (decoded_rs2[1]), .B (decoded_rs2[2]), .Y (n_988));
  NOR2X1 g181232(.A (\genblk2.pcpi_div_instr_rem ), .B
       (\genblk2.pcpi_div_instr_div ), .Y (n_987));
  NAND2XL g181233(.A (n_138), .B (n_6547), .Y (n_986));
  NOR2XL g181234(.A (pcpi_timeout), .B (instr_ecall_ebreak), .Y
       (n_985));
  OR2X1 g181235(.A (n_628), .B (n_56), .Y (n_984));
  NOR2X1 g181236(.A (mem_rdata_q[29]), .B (mem_rdata_q[28]), .Y
       (n_983));
  NOR2X1 g181237(.A (instr_srli), .B (instr_srl), .Y (n_982));
  NOR2X1 g181238(.A (is_lui_auipc_jal), .B
       (is_jalr_addi_slti_sltiu_xori_ori_andi), .Y (n_981));
  NOR2X1 g181239(.A (latched_rd[2]), .B (latched_rd[1]), .Y (n_979));
  NAND2X1 g181240(.A (n_313), .B (n_219), .Y (n_978));
  NOR2X1 g181241(.A (mem_rdata_q[26]), .B (mem_rdata_q[25]), .Y
       (n_977));
  NOR2X1 g181242(.A (latched_is_lb), .B (n_564), .Y (n_976));
  NAND2XL g181243(.A (n_6555), .B (n_543), .Y (n_975));
  NAND2X1 g181244(.A (mem_rdata_latched[1]), .B (n_345), .Y (n_974));
  NAND2X1 g181245(.A (is_lb_lh_lw_lbu_lhu), .B (n_356), .Y (n_973));
  NOR2X1 g181246(.A (n_564), .B (n_343), .Y (n_972));
  NOR2X1 g181247(.A (n_564), .B (n_311), .Y (n_971));
  AND2X1 g181248(.A (n_340), .B (cpu_state[0]), .Y (n_970));
  NOR2X1 g181249(.A (n_599), .B (n_548), .Y (n_968));
  NOR2X1 g181250(.A (n_564), .B (n_331), .Y (n_967));
  NAND2X1 g181251(.A (n_587), .B (n_580), .Y (n_966));
  NOR2X1 g181252(.A (decoded_rs1[0]), .B (decoded_rs1[2]), .Y (n_964));
  NAND2X1 g181253(.A (n_646), .B (n_593), .Y (n_963));
  NOR2BX1 g181254(.AN (is_lui_auipc_jal), .B (instr_lui), .Y (n_961));
  AND2X1 g181255(.A (decoded_rs1[2]), .B (decoded_rs1[0]), .Y (n_960));
  NOR2X1 g181256(.A (n_587), .B (n_580), .Y (n_290));
  NAND2X1 g181257(.A (decoded_rs2[4]), .B (decoded_rs2[3]), .Y (n_338));
  NOR2BX1 g181258(.AN (decoded_rs1[2]), .B (decoded_rs1[0]), .Y
       (n_957));
  AND2X2 g181260(.A (latched_store), .B (n_555), .Y (n_442));
  OR2X2 g181261(.A (\genblk2.pcpi_div_n_4742 ), .B (n_544), .Y (n_954));
  OR2X2 g181262(.A (n_602), .B (mem_done), .Y (n_953));
  OR2X4 g181263(.A (n_615), .B (n_589), .Y (n_952));
  INVX1 g181264(.A (n_883), .Y (n_884));
  INVX1 g181268(.A (n_858), .Y (n_859));
  INVX1 g181269(.A (n_848), .Y (n_847));
  INVX1 g181270(.A (n_845), .Y (n_844));
  INVX1 g181271(.A (n_843), .Y (n_842));
  AND2X1 g181281(.A (n_6782), .B (n_543), .Y (n_830));
  AND2X1 g181282(.A (n_6796), .B (n_543), .Y (n_829));
  NOR2X1 g181283(.A (cpu_state[2]), .B (cpu_state[5]), .Y (n_828));
  NAND2X1 g181284(.A (decoded_imm[29]), .B (n_537), .Y (n_827));
  AND2X1 g181285(.A (n_6757), .B (n_543), .Y (n_826));
  NOR2X1 g181286(.A (\reg_op1[16]_9653 ), .B
       (\genblk2.pcpi_div_minus_2470_59_n_481 ), .Y (n_825));
  NAND2X1 g181287(.A (mem_16bit_buffer[4]), .B (n_360), .Y (n_824));
  NAND2X1 g181288(.A (mem_16bit_buffer[2]), .B (n_360), .Y (n_823));
  AND2X1 g181289(.A (n_6762), .B (n_543), .Y (n_822));
  NAND2X1 g181290(.A (mem_16bit_buffer[7]), .B (n_360), .Y (n_821));
  NOR2X1 g181291(.A (decoder_trigger), .B (n_320), .Y (n_820));
  NAND2X1 g181292(.A (decoded_imm[27]), .B (n_537), .Y (n_819));
  AND2X1 g181293(.A (n_6755), .B (n_543), .Y (n_818));
  AND2X1 g181294(.A (n_6776), .B (n_543), .Y (n_817));
  NOR2X1 g181295(.A (\reg_op1[29]_9666 ), .B (n_721), .Y (n_816));
  AND2X1 g181296(.A (n_6785), .B (n_543), .Y (n_815));
  AND2X1 g181297(.A (n_6795), .B (n_543), .Y (n_814));
  AND2X1 g181298(.A (n_543), .B (n_6747), .Y (n_813));
  NAND2XL g181299(.A (n_6546), .B (n_6544), .Y (n_812));
  AND2X1 g181300(.A (n_6798), .B (n_543), .Y (n_811));
  NAND2X1 g181301(.A (mem_16bit_buffer[15]), .B (n_360), .Y (n_810));
  NOR2X1 g181302(.A (\reg_op2[13]_9682 ), .B (\reg_op1[13]_9650 ), .Y
       (n_809));
  AND2X1 g181303(.A (n_6760), .B (n_543), .Y (n_808));
  AND2X1 g181304(.A (n_543), .B (\genblk1.pcpi_mul_active [0]), .Y
       (n_807));
  AND2X1 g181305(.A (n_6769), .B (n_543), .Y (n_806));
  NAND2X1 g181306(.A (decoded_imm[26]), .B (n_537), .Y (n_805));
  NAND2X1 g181307(.A (n_582), .B (n_150), .Y (n_804));
  NOR2X1 g181308(.A (\reg_op2[10]_9679 ), .B (\reg_op1[10]_9647 ), .Y
       (n_803));
  AND2X1 g181309(.A (n_6772), .B (n_543), .Y (n_802));
  AND2X1 g181310(.A (n_6787), .B (n_543), .Y (n_801));
  AND2X1 g181311(.A (n_543), .B (n_6740), .Y (n_800));
  AND2X1 g181312(.A (n_543), .B (n_6745), .Y (n_799));
  NAND2X1 g181313(.A (decoded_imm[21]), .B (n_537), .Y (n_798));
  AND2X1 g181314(.A (n_6781), .B (n_543), .Y (n_797));
  AND2X1 g181315(.A (n_543), .B (n_6746), .Y (n_796));
  AND2X1 g181316(.A (n_6748), .B (n_543), .Y (n_795));
  AND2X1 g181317(.A (n_543), .B (n_6742), .Y (n_794));
  NOR2X1 g181318(.A (n_548), .B (n_356), .Y (n_793));
  NOR2X1 g181319(.A (instr_jal), .B (n_589), .Y (n_792));
  NOR2X1 g181320(.A (\reg_op2[11]_9680 ), .B (\reg_op1[11]_9648 ), .Y
       (n_791));
  AND2X1 g181321(.A (n_6797), .B (n_543), .Y (n_790));
  NOR2XL g181322(.A (last_mem_valid), .B (n_6524), .Y (n_789));
  NAND2X1 g181323(.A (mem_16bit_buffer[6]), .B (n_360), .Y (n_788));
  NAND2X1 g181324(.A (instr_sltiu), .B (n_537), .Y (n_787));
  NAND2X1 g181325(.A (mem_16bit_buffer[9]), .B (n_360), .Y (n_786));
  NOR2X1 g181326(.A (\reg_op2[18]_9687 ), .B (\reg_op1[18]_9655 ), .Y
       (n_785));
  AND2X1 g181327(.A (n_6792), .B (n_543), .Y (n_784));
  AND2X1 g181328(.A (n_6783), .B (n_543), .Y (n_783));
  AND2X1 g181329(.A (n_6766), .B (n_543), .Y (n_782));
  NAND2X1 g181330(.A (instr_sub), .B (n_537), .Y (n_781));
  NAND2X1 g181331(.A (decoded_rs2[1]), .B (decoded_rs2[2]), .Y (n_885));
  NOR2X1 g181333(.A (\reg_op1[8]_9645 ), .B
       (\genblk2.pcpi_div_minus_2470_59_n_492 ), .Y (n_883));
  NOR2X1 g181334(.A (decoded_rs2[1]), .B (n_651), .Y (n_882));
  NOR2X1 g181335(.A (n_595), .B (n_219), .Y (n_881));
  NAND2X1 g181336(.A (decoded_rs2[1]), .B (n_651), .Y (n_880));
  NOR2X1 g181337(.A (\reg_op1[9]_9646 ), .B (n_714), .Y (n_879));
  NOR2X1 g181338(.A (reg_op1[0]), .B (n_630), .Y (n_878));
  NAND2X1 g181339(.A (mem_rdata_q[14]), .B (mem_rdata_q[13]), .Y
       (n_877));
  NAND2XL g181340(.A (n_6550), .B (n_6549), .Y (n_876));
  NOR2X1 g181342(.A (cpu_state[6]), .B (cpu_state[3]), .Y (n_779));
  NAND2X1 g181343(.A (is_beq_bne_blt_bge_bltu_bgeu), .B (n_538), .Y
       (n_875));
  NAND2X1 g181344(.A (mem_rdata_q[14]), .B (n_640), .Y (n_874));
  NOR2X1 g181345(.A (\reg_op1[6]_9643 ), .B
       (\genblk2.pcpi_div_minus_2470_59_n_474 ), .Y (n_873));
  NAND2X1 g181347(.A (\reg_op1[18]_9655 ), .B
       (\genblk2.pcpi_div_minus_2470_59_n_485 ), .Y (n_871));
  NAND2X1 g181348(.A (\reg_op1[6]_9643 ), .B
       (\genblk2.pcpi_div_minus_2470_59_n_474 ), .Y (n_870));
  NAND2X1 g181349(.A (\reg_op1[12]_9649 ), .B
       (\genblk2.pcpi_div_minus_2470_59_n_498 ), .Y (n_869));
  NAND2X1 g181350(.A (\reg_op2[31]_9700 ), .B (n_627), .Y (n_868));
  NAND2X1 g181351(.A (\reg_op1[14]_9651 ), .B
       (\genblk2.pcpi_div_minus_2470_59_n_499 ), .Y (n_867));
  NOR2X1 g181352(.A (\reg_op2[31]_9700 ), .B (n_627), .Y (n_866));
  NAND2X1 g181353(.A (\reg_op1[13]_9650 ), .B (n_572), .Y (n_865));
  NAND2X1 g181355(.A (\reg_op2[7]_9676 ), .B (n_744), .Y (n_863));
  NAND2X1 g181356(.A (\reg_op2[14]_9683 ), .B (n_624), .Y (n_862));
  NAND2X1 g181357(.A (\reg_op1[11]_9648 ), .B (n_751), .Y (n_861));
  NAND2X1 g181359(.A (\reg_op1[10]_9647 ), .B
       (\genblk2.pcpi_div_minus_2470_59_n_502 ), .Y (n_860));
  NAND2X1 g181360(.A (\reg_op1[15]_9652 ), .B (n_635), .Y (n_858));
  NAND2X1 g181361(.A (\reg_op2[18]_9687 ), .B (n_625), .Y (n_857));
  NOR2X1 g181362(.A (\reg_op2[7]_9676 ), .B (n_744), .Y (n_856));
  NAND2X1 g181363(.A (\reg_op2[15]_9684 ), .B (n_619), .Y (n_855));
  NAND2X1 g181364(.A (\reg_op1[31]_9668 ), .B (cpu_state[2]), .Y
       (n_854));
  NAND2X1 g181365(.A (mem_rdata_q[13]), .B (n_641), .Y (n_853));
  NAND2X1 g181366(.A (n_564), .B (n_611), .Y (n_852));
  NAND2X1 g181367(.A (is_sb_sh_sw), .B (n_538), .Y (n_851));
  NAND2X1 g181369(.A (n_543), .B (mem_done), .Y (n_850));
  NOR2X1 g181370(.A (is_beq_bne_blt_bge_bltu_bgeu), .B (n_613), .Y
       (n_849));
  NAND2X1 g181371(.A (n_587), .B (latched_rd[3]), .Y (n_848));
  NOR2BX1 g181372(.AN (decoded_rs1[0]), .B (decoded_rs1[2]), .Y
       (n_846));
  NOR2X1 g181373(.A (n_587), .B (latched_rd[3]), .Y (n_845));
  NAND2X1 g181374(.A (decoded_rs2[3]), .B (n_593), .Y (n_843));
  NAND2X1 g181375(.A (decoded_rs2[4]), .B (n_646), .Y (n_289));
  NOR2X1 g181376(.A (n_5693), .B (n_544), .Y (n_545));
  AND2X1 g181377(.A (n_446), .B (mem_la_secondword), .Y (n_839));
  NOR2X1 g181378(.A (n_562), .B (n_446), .Y (n_505));
  AND2X1 g181379(.A (n_538), .B (instr_jal), .Y (n_441));
  AND2X2 g181382(.A (n_615), .B (n_543), .Y (n_427));
  OR2X2 g181383(.A (cpu_state[1]), .B (cpu_state[0]), .Y (n_833));
  OR2X2 g181384(.A (n_548), .B (n_544), .Y (n_832));
  NAND2X1 g181385(.A (cpu_state[6]), .B (n_543), .Y (n_324));
  INVXL g181386(.A (n_6551), .Y (n_778));
  INVX1 g181388(.A (decoded_rd[3]), .Y (n_777));
  INVX1 g181390(.A (decoded_imm_j[10]), .Y (n_776));
  INVX1 g181404(.A (decoded_imm_j[16]), .Y (n_775));
  INVX1 g181409(.A (decoded_imm_j[15]), .Y (n_774));
  INVX1 g181438(.A (pcpi_mul_wr), .Y (n_773));
  INVX1 g181477(.A (decoded_imm_j[7]), .Y (n_772));
  INVX1 g181489(.A (decoded_imm_j[11]), .Y (n_771));
  INVX1 g181509(.A (pcpi_timeout_counter[0]), .Y (n_770));
  INVX1 g181518(.A (decoded_imm_j[6]), .Y (n_769));
  INVX1 g181521(.A (decoded_imm[5]), .Y (n_768));
  INVX1 g181525(.A (is_sll_srl_sra), .Y (n_767));
  INVX1 g181549(.A (instr_srai), .Y (n_766));
  INVX1 g181570(.A (decoded_imm[7]), .Y (n_765));
  INVX1 g181581(.A (mem_state[0]), .Y (n_764));
  INVX1 g181596(.A (mem_rdata_q[2]), .Y (n_763));
  INVX1 g181598(.A (mem_rdata_q[16]), .Y (n_762));
  INVX1 g181607(.A (cpu_state[1]), .Y (n_761));
  INVX1 g181612(.A (\reg_op2[27]_9696 ), .Y (n_760));
  INVX1 g181627(.A (mem_rdata_q[0]), .Y (n_759));
  INVX1 g181633(.A (\reg_op2[20]_9689 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_500 ));
  INVX1 g181642(.A (\reg_op2[2]_9671 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_487 ));
  INVX1 g181654(.A (\reg_op2[26]_9695 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_488 ));
  INVX1 g181671(.A (mem_rdata_q[29]), .Y (n_752));
  INVX1 g181680(.A (\reg_op2[11]_9680 ), .Y (n_751));
  INVX1 g181697(.A (\reg_op1[21]_9658 ), .Y (n_637));
  INVX1 g181702(.A (\reg_op2[14]_9683 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_499 ));
  INVX1 g181711(.A (\reg_op2[18]_9687 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_485 ));
  INVX1 g181723(.A (\reg_op2[15]_9684 ), .Y (n_635));
  INVX1 g181732(.A (\reg_op2[10]_9679 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_502 ));
  INVX1 g181742(.A (\reg_op1[19]_9656 ), .Y (n_747));
  INVX1 g181769(.A (\reg_op2[8]_9677 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_492 ));
  INVX1 g181772(.A (\reg_op2[7]_9676 ), .Y (n_746));
  INVX1 g181803(.A (n_46), .Y (n_745));
  INVX1 g181816(.A (\reg_op2[0]_9669 ), .Y (n_630));
  INVX1 g181829(.A (\reg_op2[1]_9670 ), .Y (n_629));
  INVX1 g181848(.A (reg_op1[0]), .Y (n_628));
  INVX1 g181863(.A (\reg_op1[31]_9668 ), .Y (n_627));
  INVX1 g181884(.A (\reg_op1[18]_9655 ), .Y (n_625));
  INVX1 g181905(.A (\reg_op1[14]_9651 ), .Y (n_624));
  INVX1 g181921(.A (\reg_op1[7]_9644 ), .Y (n_744));
  INVX1 g181953(.A (\reg_op1[15]_9652 ), .Y (n_619));
  INVX1 g181990(.A (decoded_rd[2]), .Y (n_740));
  INVX1 g181991(.A (n_42), .Y (n_739));
  INVX1 g181995(.A (decoded_rd[1]), .Y (n_736));
  INVX1 g182011(.A (decoded_imm_j[19]), .Y (n_735));
  INVX1 g182068(.A (\genblk2.pcpi_div_quotient_msk [0]), .Y (n_734));
  INVX1 g182070(.A (decoded_imm_j[5]), .Y (n_733));
  INVX1 g182074(.A (decoded_imm[10]), .Y (n_732));
  INVX1 g182105(.A (decoded_imm_j[17]), .Y (n_731));
  INVX1 g182166(.A (decoded_imm[6]), .Y (n_730));
  INVX1 g182184(.A (is_alu_reg_reg), .Y (n_729));
  INVX1 g182193(.A (mem_rdata_q[17]), .Y (n_728));
  INVX1 g182205(.A (mem_rdata_q[28]), .Y (n_727));
  INVX1 g182211(.A (decoder_trigger), .Y (n_589));
  INVX1 g182214(.A (\reg_op2[17]_9686 ), .Y (n_726));
  INVX1 g182226(.A (\reg_op2[28]_9697 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_479 ));
  INVX1 g182236(.A (instr_jalr), .Y (n_723));
  INVX1 g182240(.A (\reg_op2[25]_9694 ), .Y (n_722));
  INVX1 g182247(.A (\reg_op2[29]_9698 ), .Y (n_721));
  INVX1 g182260(.A (\reg_op2[16]_9685 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_481 ));
  INVX1 g182265(.A (\reg_op2[24]_9693 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_483 ));
  INVX1 g182298(.A (\reg_op1[3]_9640 ), .Y (n_578));
  INVX1 g182306(.A (\reg_op1[2]_9639 ), .Y (n_577));
  INVX1 g182312(.A (\reg_op1[22]_9659 ), .Y (n_576));
  INVX1 g182326(.A (\reg_op2[12]_9681 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_498 ));
  INVX1 g182353(.A (\reg_op2[31]_9700 ), .Y (n_573));
  INVX1 g182358(.A (\reg_op2[13]_9682 ), .Y (n_572));
  INVX1 g182390(.A (\reg_op2[6]_9675 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_474 ));
  INVX1 g182402(.A (\reg_op2[9]_9678 ), .Y (n_714));
  INVX1 g182440(.A (n_113), .Y (n_712));
  INVX1 g182485(.A (\reg_op1[1]_9638 ), .Y (n_565));
  INVX1 g182501(.A (cpu_state[0]), .Y (n_564));
  INVX1 g182509(.A (mem_la_secondword), .Y (n_562));
  INVX1 g182539(.A (instr_rdinstr), .Y (n_709));
  INVX1 g182557(.A (instr_rdcycle), .Y (n_707));
  INVX1 g182571(.A (latched_branch), .Y (n_555));
  DFFX1 clear_prefetched_high_word_q_reg(.CK (clk), .D (n_1167), .Q
       (clear_prefetched_high_word_q), .QN (n_654));
  DFFX2 \cpu_state_reg[2] (.CK (clk), .D (n_5067), .Q (cpu_state[2]),
       .QN (n_611));
  DFFX2 \cpu_state_reg[3] (.CK (clk), .D (n_5069), .Q (cpu_state[3]),
       .QN (n_613));
  DFFX1 \cpu_state_reg[6] (.CK (clk), .D (n_5121), .Q (cpu_state[6]),
       .QN (n_615));
  DFFX1 \cpuregs_reg[3][19] (.CK (clk), .D (n_4196), .Q
       (\cpuregs[3] [19]), .QN (n_604));
  DFFX1 \cpuregs_reg[3][21] (.CK (clk), .D (n_4203), .Q
       (\cpuregs[3] [21]), .QN (n_655));
  DFFX1 \cpuregs_reg[3][22] (.CK (clk), .D (n_4206), .Q
       (\cpuregs[3] [22]), .QN (n_606));
  DFFX1 \decoded_imm_reg[0] (.CK (clk), .D (n_2179), .Q
       (decoded_imm[0]), .QN (n_605));
  DFFX1 \decoded_rs1_reg[4] (.CK (clk), .D (n_4734), .Q
       (decoded_rs1[4]), .QN (n_574));
  DFFX1 \decoded_rs2_reg[0] (.CK (clk), .D (n_4847), .Q
       (decoded_rs2[0]), .QN (n_633));
  DFFX1 \decoded_rs2_reg[2] (.CK (clk), .D (n_4848), .Q
       (decoded_rs2[2]), .QN (n_651));
  DFFX1 \decoded_rs2_reg[3] (.CK (clk), .D (n_4758), .Q
       (decoded_rs2[3]), .QN (n_646));
  DFFX1 \decoded_rs2_reg[4] (.CK (clk), .D (n_4532), .Q
       (decoded_rs2[4]), .QN (n_593));
  DFFX1 instr_jal_reg(.CK (clk), .D (n_3017), .Q (instr_jal), .QN
       (n_652));
  DFFX1 is_alu_reg_imm_reg(.CK (clk), .D (n_4846), .Q (is_alu_reg_imm),
       .QN (n_622));
  DFFX1 is_slli_srli_srai_reg(.CK (clk), .D (n_3018), .Q
       (is_slli_srli_srai), .QN (n_599));
  DFFX1 \latched_rd_reg[1] (.CK (clk), .D (n_1746), .Q (latched_rd[1]),
       .QN (n_592));
  DFFX1 \latched_rd_reg[2] (.CK (clk), .D (n_1742), .Q (latched_rd[2]),
       .QN (n_638));
  DFFX1 \latched_rd_reg[3] (.CK (clk), .D (n_1745), .Q (latched_rd[3]),
       .QN (n_580));
  DFFX1 \latched_rd_reg[4] (.CK (clk), .D (n_1744), .Q (latched_rd[4]),
       .QN (n_587));
  DFFX1 mem_do_prefetch_reg(.CK (clk), .D (n_2305), .Q
       (mem_do_prefetch), .QN (n_595));
  DFFX1 mem_do_rdata_reg(.CK (clk), .D (n_2418), .Q (mem_do_rdata), .QN
       (n_582));
  DFFX1 mem_do_rinst_reg(.CK (clk), .D (n_5523), .Q (mem_do_rinst), .QN
       (n_602));
  DFFX1 \mem_rdata_q_reg[4] (.CK (clk), .D (n_2342), .Q
       (mem_rdata_q[4]), .QN (n_594));
  DFFX1 \mem_rdata_q_reg[5] (.CK (clk), .D (n_2341), .Q
       (mem_rdata_q[5]), .QN (n_649));
  DFFX1 \mem_rdata_q_reg[6] (.CK (clk), .D (n_2340), .Q
       (mem_rdata_q[6]), .QN (n_586));
  DFFX1 \mem_rdata_q_reg[7] (.CK (clk), .D (n_4855), .Q
       (mem_rdata_q[7]), .QN (n_643));
  DFFX1 \mem_rdata_q_reg[8] (.CK (clk), .D (n_4853), .Q
       (mem_rdata_q[8]), .QN (n_647));
  DFFX1 \mem_rdata_q_reg[9] (.CK (clk), .D (n_4096), .Q
       (mem_rdata_q[9]), .QN (n_650));
  DFFX1 \mem_rdata_q_reg[12] (.CK (clk), .D (n_5178), .Q
       (mem_rdata_q[12]), .QN (n_616));
  DFFX1 \mem_rdata_q_reg[13] (.CK (clk), .D (n_5235), .Q
       (mem_rdata_q[13]), .QN (n_640));
  DFFX1 \mem_rdata_q_reg[14] (.CK (clk), .D (n_5125), .Q
       (mem_rdata_q[14]), .QN (n_641));
  DFFX1 \mem_rdata_q_reg[15] (.CK (clk), .D (n_4714), .Q
       (mem_rdata_q[15]), .QN (n_583));
  DFFX1 \mem_rdata_q_reg[18] (.CK (clk), .D (n_4733), .Q
       (mem_rdata_q[18]), .QN (n_596));
  DFFX1 \mem_rdata_q_reg[19] (.CK (clk), .D (n_4735), .Q
       (mem_rdata_q[19]), .QN (n_597));
  DFFX1 \mem_rdata_q_reg[20] (.CK (clk), .D (n_5118), .Q
       (mem_rdata_q[20]), .QN (n_588));
  DFFX1 \mem_rdata_q_reg[21] (.CK (clk), .D (n_5120), .Q
       (mem_rdata_q[21]), .QN (n_644));
  DFFX1 \mem_rdata_q_reg[22] (.CK (clk), .D (n_5122), .Q
       (mem_rdata_q[22]), .QN (n_581));
  DFFX1 \mem_rdata_q_reg[23] (.CK (clk), .D (n_5117), .Q
       (mem_rdata_q[23]), .QN (n_639));
  DFFX1 \mem_rdata_q_reg[24] (.CK (clk), .D (n_5123), .Q
       (mem_rdata_q[24]), .QN (n_590));
  DFFX1 \mem_rdata_q_reg[25] (.CK (clk), .D (n_5229), .Q
       (mem_rdata_q[25]), .QN (n_648));
  DFFX1 \mem_rdata_q_reg[26] (.CK (clk), .D (n_5170), .Q
       (mem_rdata_q[26]), .QN (n_591));
  DFFX1 \mem_rdata_q_reg[27] (.CK (clk), .D (n_5169), .Q
       (mem_rdata_q[27]), .QN (n_642));
  DFFX1 \mem_rdata_q_reg[30] (.CK (clk), .D (n_5200), .Q
       (mem_rdata_q[30]), .QN (n_579));
  DFFX1 \mem_rdata_q_reg[31] (.CK (clk), .D (n_5151), .Q
       (mem_rdata_q[31]), .QN (n_636));
  DFFX1 \mem_state_reg[1] (.CK (clk), .D (n_3176), .Q (mem_state[1]),
       .QN (n_603));
  INVX1 drc_bufs183002(.A (n_550), .Y (n_677));
  INVX1 drc_bufs183025(.A (n_545), .Y (n_664));
  INVX3 drc_bufs183055(.A (n_952), .Y (n_666));
  INVX1 drc_bufs183083(.A (n_954), .Y (n_668));
  INVX1 drc_bufs183091(.A (n_953), .Y (n_667));
  INVX1 drc_bufs183097(.A (n_13034), .Y (n_540));
  INVX3 drc_bufs183113(.A (n_538), .Y (n_537));
  INVX1 drc_bufs183135(.A (n_832), .Y (n_659));
  INVX1 drc_bufs183263(.A (n_3219), .Y (n_697));
  INVX1 drc_bufs183282(.A (n_505), .Y (n_663));
  INVX1 drc_bufs183391(.A (n_504), .Y (n_680));
  INVX2 drc_bufs183639(.A (n_445), .Y (n_446));
  INVX2 drc_bufs183640(.A (mem_xfer), .Y (n_445));
  INVX1 drc_bufs183662(.A (n_441), .Y (n_662));
  INVX1 drc_bufs183673(.A (n_440), .Y (n_681));
  INVX1 drc_bufs183678(.A (n_439), .Y (n_688));
  INVX1 drc_bufs183682(.A (n_438), .Y (n_685));
  INVX1 drc_bufs183686(.A (n_437), .Y (n_682));
  INVX1 drc_bufs183719(.A (n_432), .Y (n_704));
  INVX1 drc_bufs183772(.A (n_33), .Y (n_419));
  INVX1 drc_bufs184036(.A (n_356), .Y (n_645));
  INVX1 drc_bufs184057(.A (n_32), .Y (n_349));
  INVX1 drc_bufs184063(.A (n_348), .Y (n_702));
  INVX1 drc_bufs184067(.A (n_347), .Y (n_695));
  INVX1 drc_bufs184071(.A (mem_rdata_latched[0]), .Y (n_345));
  INVX1 drc_bufs184080(.A (n_344), .Y (n_691));
  INVX1 drc_bufs184083(.A (n_343), .Y (n_607));
  INVX1 drc_bufs184087(.A (n_342), .Y (n_673));
  INVX1 drc_bufs184093(.A (n_341), .Y (n_703));
  INVX1 drc_bufs184173(.A (n_335), .Y (n_674));
  INVX1 drc_bufs184194(.A (n_334), .Y (n_679));
  INVX1 drc_bufs184211(.A (n_332), .Y (n_678));
  INVX1 drc_bufs184223(.A (n_327), .Y (n_687));
  INVX1 drc_bufs184227(.A (n_326), .Y (n_689));
  INVX1 drc_bufs184231(.A (n_325), .Y (n_690));
  INVX2 drc_bufs184235(.A (n_324), .Y (n_658));
  INVX1 drc_bufs184247(.A (n_693), .Y (n_321));
  INVX1 drc_bufs184248(.A (n_2489), .Y (n_693));
  INVX1 drc_bufs184276(.A (n_30), .Y (n_314));
  INVX1 drc_bufs184288(.A (n_29), .Y (n_310));
  INVX1 drc_bufs184292(.A (n_28), .Y (n_309));
  INVX1 drc_bufs184298(.A (n_308), .Y (n_696));
  INVX1 drc_bufs184300(.A (n_27), .Y (n_307));
  INVX1 drc_bufs184304(.A (n_26), .Y (n_306));
  INVX1 drc_bufs184312(.A (n_25), .Y (n_303));
  INVX1 drc_bufs184316(.A (n_24), .Y (n_302));
  INVX1 drc_bufs184322(.A (n_301), .Y (n_705));
  INVX1 drc_bufs184324(.A (n_23), .Y (n_300));
  INVX1 drc_bufs184332(.A (n_22), .Y (n_297));
  INVX1 drc_bufs184346(.A (n_294), .Y (n_706));
  INVX1 drc_bufs184362(.A (n_2435), .Y (n_692));
  INVX1 drc_bufs184366(.A (n_290), .Y (n_671));
  INVX1 drc_bufs184382(.A (n_1310), .Y (n_672));
  INVX1 drc_bufs184385(.A (n_289), .Y (n_665));
  INVX1 drc_bufs184389(.A (n_1319), .Y (n_675));
  INVX1 drc_bufs184393(.A (n_1322), .Y (n_676));
  INVX1 drc_bufs184405(.A (n_2137), .Y (n_683));
  INVX1 drc_bufs184409(.A (n_2140), .Y (n_686));
  BUFX20 fopt184451(.A (n_5655), .Y (mem_wdata[25]));
  BUFX20 fopt184453(.A (n_5651), .Y (mem_wdata[21]));
  BUFX20 fopt184455(.A (n_5641), .Y (mem_wdata[11]));
  BUFX20 fopt184457(.A (n_5643), .Y (mem_wdata[13]));
  BUFX20 fopt184459(.A (n_5659), .Y (mem_wdata[29]));
  BUFX20 fopt184461(.A (n_5693), .Y (trap));
  BUFX20 fopt184463(.A (n_5691), .Y (mem_addr[31]));
  BUFX20 fopt184465(.A (n_5638), .Y (mem_wdata[8]));
  BUFX20 fopt184467(.A (n_5637), .Y (mem_wdata[7]));
  BUFX20 fopt184469(.A (n_5639), .Y (mem_wdata[9]));
  BUFX20 fopt184471(.A (n_5635), .Y (mem_wdata[5]));
  BUFX20 fopt184473(.A (n_5634), .Y (mem_wdata[4]));
  BUFX20 fopt184475(.A (n_5667), .Y (mem_addr[7]));
  BUFX20 fopt184477(.A (n_5633), .Y (mem_wdata[3]));
  BUFX20 fopt184479(.A (n_5636), .Y (mem_wdata[6]));
  BUFX20 fopt184481(.A (n_5631), .Y (mem_wdata[1]));
  BUFX20 fopt184483(.A (n_5671), .Y (mem_addr[11]));
  BUFX20 fopt184485(.A (n_5640), .Y (mem_wdata[10]));
  BUFX20 fopt184487(.A (n_5630), .Y (mem_wdata[0]));
  BUFX20 fopt184489(.A (n_5629), .Y (mem_wstrb[3]));
  BUFX20 fopt184491(.A (n_5675), .Y (mem_addr[15]));
  BUFX20 fopt184493(.A (n_5627), .Y (mem_wstrb[1]));
  BUFX20 fopt184495(.A (n_5632), .Y (mem_wdata[2]));
  BUFX20 fopt184497(.A (n_5628), .Y (mem_wstrb[2]));
  BUFX20 fopt184499(.A (n_5626), .Y (mem_wstrb[0]));
  BUFX20 fopt184501(.A (n_5692), .Y (mem_instr));
  BUFX20 fopt184503(.A (n_5690), .Y (mem_addr[30]));
  BUFX20 fopt184505(.A (n_5609), .Y (pcpi_insn[24]));
  BUFX20 fopt184507(.A (n_5683), .Y (mem_addr[23]));
  BUFX20 fopt184509(.A (n_5689), .Y (mem_addr[29]));
  BUFX20 fopt184511(.A (n_5608), .Y (pcpi_insn[23]));
  BUFX20 fopt184513(.A (n_5607), .Y (pcpi_insn[22]));
  BUFX20 fopt184515(.A (n_5592), .Y (pcpi_insn[7]));
  BUFX20 fopt184517(.A (n_5606), .Y (pcpi_insn[21]));
  BUFX20 fopt184519(.A (n_5605), .Y (pcpi_insn[20]));
  BUFX20 fopt184521(.A (n_5604), .Y (pcpi_insn[19]));
  BUFX20 fopt184523(.A (n_5603), .Y (pcpi_insn[18]));
  BUFX20 fopt184525(.A (n_5602), .Y (pcpi_insn[17]));
  BUFX20 fopt184527(.A (n_5601), .Y (pcpi_insn[16]));
  BUFX20 fopt184529(.A (n_5688), .Y (mem_addr[28]));
  BUFX20 fopt184531(.A (n_5600), .Y (pcpi_insn[15]));
  BUFX20 fopt184533(.A (n_5596), .Y (pcpi_insn[11]));
  BUFX20 fopt184535(.A (n_5595), .Y (pcpi_insn[10]));
  BUFX20 fopt184537(.A (n_5594), .Y (pcpi_insn[9]));
  BUFX20 fopt184539(.A (n_5687), .Y (mem_addr[27]));
  BUFX20 fopt184541(.A (n_5593), .Y (pcpi_insn[8]));
  BUFX20 fopt184543(.A (n_5686), .Y (mem_addr[26]));
  BUFX20 fopt184545(.A (n_5685), .Y (mem_addr[25]));
  BUFX20 fopt184547(.A (n_5684), .Y (mem_addr[24]));
  BUFX20 fopt184549(.A (n_5681), .Y (mem_addr[21]));
  BUFX20 fopt184551(.A (n_5680), .Y (mem_addr[20]));
  BUFX20 fopt184553(.A (n_5679), .Y (mem_addr[19]));
  BUFX20 fopt184555(.A (n_5678), .Y (mem_addr[18]));
  BUFX20 fopt184557(.A (n_5677), .Y (mem_addr[17]));
  BUFX20 fopt184559(.A (n_5676), .Y (mem_addr[16]));
  BUFX20 fopt184561(.A (n_5674), .Y (mem_addr[14]));
  BUFX20 fopt184563(.A (n_5673), .Y (mem_addr[13]));
  BUFX20 fopt184565(.A (n_5672), .Y (mem_addr[12]));
  BUFX20 fopt184567(.A (n_5670), .Y (mem_addr[10]));
  BUFX20 fopt184569(.A (n_5669), .Y (mem_addr[9]));
  BUFX20 fopt184571(.A (n_5668), .Y (mem_addr[8]));
  BUFX20 fopt184573(.A (n_5666), .Y (mem_addr[6]));
  BUFX20 fopt184575(.A (n_5665), .Y (mem_addr[5]));
  BUFX20 fopt184577(.A (n_5664), .Y (mem_addr[4]));
  BUFX20 fopt184579(.A (n_5663), .Y (mem_addr[3]));
  BUFX20 fopt184581(.A (n_5662), .Y (mem_addr[2]));
  BUFX20 fopt184583(.A (n_5661), .Y (mem_wdata[31]));
  BUFX20 fopt184585(.A (n_5660), .Y (mem_wdata[30]));
  BUFX20 fopt184587(.A (n_5658), .Y (mem_wdata[28]));
  BUFX20 fopt184589(.A (n_5657), .Y (mem_wdata[27]));
  BUFX20 fopt184591(.A (n_5656), .Y (mem_wdata[26]));
  BUFX20 fopt184593(.A (n_5654), .Y (mem_wdata[24]));
  BUFX20 fopt184595(.A (n_5653), .Y (mem_wdata[23]));
  BUFX20 fopt184597(.A (n_5652), .Y (mem_wdata[22]));
  BUFX20 fopt184599(.A (n_5648), .Y (mem_wdata[18]));
  BUFX20 fopt184601(.A (n_5647), .Y (mem_wdata[17]));
  BUFX20 fopt184603(.A (n_5646), .Y (mem_wdata[16]));
  BUFX20 fopt184605(.A (n_5645), .Y (mem_wdata[15]));
  BUFX20 fopt184607(.A (n_5644), .Y (mem_wdata[14]));
  BUFX20 fopt184609(.A (n_5682), .Y (mem_addr[22]));
  BUFX20 fopt184611(.A (n_5649), .Y (mem_wdata[19]));
  BUFX20 fopt184613(.A (n_5642), .Y (mem_wdata[12]));
  BUFX20 fopt184615(.A (n_5650), .Y (mem_wdata[20]));
  INVX3 drc_bufs184625(.A (n_544), .Y (n_543));
  CLKINVX6 drc_bufs184629(.A (resetn), .Y (n_544));
  INVX1 drc_bufs184665(.A (n_279), .Y (n_278));
  INVX1 drc_bufs184712(.A (mem_rdata[25]), .Y (n_653));
  INVX1 drc_bufs184716(.A (mem_rdata[15]), .Y (n_600));
  INVX1 drc_bufs184789(.A (mem_rdata[9]), .Y (n_601));
  INVX1 drc_bufs184793(.A (mem_rdata[31]), .Y (n_598));
  INVX1 drc_bufs184801(.A (mem_done), .Y (n_219));
  INVX1 drc_bufs185007(.A (mem_rdata[7]), .Y (n_656));
  INVX1 drc_bufs185204(.A (\genblk2.pcpi_div_n_314 ), .Y (n_609));
  INVX3 drc_bufs185674(.A (n_40), .Y (n_39));
  AND2X1 g91915(.A (n_344), .B (n_1621), .Y (n_38));
  OAI2BB1X2 g186344(.A0N (n_1543), .A1N (n_1951), .B0 (cpu_state[0]),
       .Y (n_37));
  AOI21X1 g186345(.A0 (decoded_imm_j[20]), .A1 (n_441), .B0 (n_2162),
       .Y (n_36));
  NAND3X1 g186346(.A (n_445), .B (n_2510), .C (n_2604), .Y (n_35));
  OAI31X1 g186347(.A0 (instr_jalr), .A1 (is_alu_reg_imm), .A2
       (is_lb_lh_lw_lbu_lhu), .B0 (n_538), .Y (n_34));
  OR3X1 g186348(.A (mem_rdata_latched[1]), .B (mem_rdata_latched[0]),
       .C (n_335), .Y (n_33));
  AND4X1 g186349(.A (n_2822), .B (n_667), .C (n_342), .D (n_3015), .Y
       (n_32));
  AND4X1 g186350(.A (n_317), .B (n_2433), .C (n_2600), .D (n_429), .Y
       (n_31));
  AND4X1 g186351(.A (mem_state[0]), .B (n_582), .C (n_545), .D
       (n_2430), .Y (n_30));
  AND4X1 g186352(.A (n_2050), .B (n_2070), .C (n_2310), .D (n_3166), .Y
       (n_29));
  AND4X1 g186353(.A (n_2051), .B (n_2041), .C (n_2311), .D (n_3167), .Y
       (n_28));
  OR3X1 g186354(.A (pcpi_div_wait), .B (pcpi_wait), .C (n_989), .Y
       (n_27));
  AND4X1 g186355(.A (mem_rdata_q[31]), .B (mem_rdata_q[30]), .C
       (n_1326), .D (n_3430), .Y (n_26));
  AND4X1 g186356(.A (n_1357), .B (n_2165), .C (n_2484), .D (n_1361), .Y
       (n_25));
  AND4X1 g186357(.A (n_2140), .B (n_683), .C (n_682), .D (n_673), .Y
       (n_24));
  AND4X1 g186358(.A (n_2018), .B (n_2068), .C (n_2066), .D (n_3193), .Y
       (n_23));
  AND4X1 g186359(.A (n_288), .B (n_6527), .C (n_40), .D (n_917), .Y
       (n_22));
  NAND2BX1 g186360(.AN (latched_rd[2]), .B (n_3004), .Y (n_21));
  NAND2BX1 g186361(.AN (n_3002), .B (decoded_rs1[1]), .Y (n_20));
  NOR2BX1 g186362(.AN (n_3001), .B (n_638), .Y (n_19));
  NOR2BX1 g186363(.AN (n_2607), .B (n_2423), .Y (n_18));
  NOR2X4 g186364(.A (n_1331), .B (n_2598), .Y (n_506));
  NOR2BX1 g186365(.AN (n_2440), .B (n_1329), .Y (n_17));
  NAND2BX1 g186366(.AN (n_2338), .B (reg_sh[4]), .Y (n_16));
  NAND2BX1 g186367(.AN (n_2320), .B (n_690), .Y (n_15));
  NOR2BX1 g186368(.AN (n_1620), .B (n_2438), .Y (n_14));
  NOR2BX1 g186369(.AN (n_1619), .B (n_2434), .Y (n_13));
  NOR2BX4 g186370(.AN (n_1602), .B (n_691), .Y (n_12));
  NOR2BX1 g186371(.AN (n_1355), .B (cpu_state[7]), .Y (n_11));
  NOR2BX1 g186372(.AN (n_1335), .B (n_289), .Y (n_10));
  NOR2BX1 g186373(.AN (n_8), .B (n_338), .Y (n_9));
  NOR2BX1 g186374(.AN (n_882), .B (decoded_rs2[0]), .Y (n_8));
  NAND2BX1 g186375(.AN (n_880), .B (decoded_rs2[0]), .Y (n_7));
  NAND2BX1 g186376(.AN (n_879), .B (n_1350), .Y (n_6));
  NAND2BX1 g186377(.AN (\reg_op1[11]_9648 ), .B (\reg_op2[11]_9680 ),
       .Y (n_5));
  NOR2BX1 g186378(.AN (\reg_op1[26]_9663 ), .B (n_1943), .Y (n_4));
  NAND2BX1 g186379(.AN (\reg_op1[10]_9647 ), .B (\reg_op2[10]_9679 ),
       .Y (n_3));
  NAND2BX1 g186380(.AN (n_833), .B (n_548), .Y (n_2));
  AO21X1 g186381(.A0 (n_2433), .A1 (n_2995), .B0 (n_31), .Y (n_1));
  NOR2BX1 g186382(.AN (n_608), .B (n_739), .Y (n_0));
  XNOR2X1 inc_add_1559_34_g848(.A (count_instr[63]), .B
       (inc_add_1559_34_n_445), .Y (n_6992));
  OA21X1 inc_add_1559_34_g849(.A0 (count_instr[62]), .A1
       (inc_add_1559_34_n_450), .B0 (inc_add_1559_34_n_445), .Y
       (n_6993));
  NAND2X1 inc_add_1559_34_g850(.A (count_instr[62]), .B
       (inc_add_1559_34_n_450), .Y (inc_add_1559_34_n_445));
  XNOR2X1 inc_add_1559_34_g851(.A (count_instr[61]), .B
       (inc_add_1559_34_n_455), .Y (n_6994));
  NOR2BX1 inc_add_1559_34_g852(.AN (count_instr[61]), .B
       (inc_add_1559_34_n_455), .Y (inc_add_1559_34_n_450));
  OA21X1 inc_add_1559_34_g853(.A0 (count_instr[60]), .A1
       (inc_add_1559_34_n_460), .B0 (inc_add_1559_34_n_455), .Y
       (n_6995));
  NAND2X1 inc_add_1559_34_g854(.A (count_instr[60]), .B
       (inc_add_1559_34_n_460), .Y (inc_add_1559_34_n_455));
  XNOR2X1 inc_add_1559_34_g855(.A (count_instr[59]), .B
       (inc_add_1559_34_n_465), .Y (n_6996));
  NOR2BX1 inc_add_1559_34_g856(.AN (count_instr[59]), .B
       (inc_add_1559_34_n_465), .Y (inc_add_1559_34_n_460));
  OA21X1 inc_add_1559_34_g857(.A0 (count_instr[58]), .A1
       (inc_add_1559_34_n_470), .B0 (inc_add_1559_34_n_465), .Y
       (n_6997));
  NAND2X1 inc_add_1559_34_g858(.A (count_instr[58]), .B
       (inc_add_1559_34_n_470), .Y (inc_add_1559_34_n_465));
  AOI2BB1X1 inc_add_1559_34_g859(.A0N (count_instr[57]), .A1N
       (inc_add_1559_34_n_475), .B0 (inc_add_1559_34_n_470), .Y
       (n_6998));
  AND2X1 inc_add_1559_34_g860(.A (inc_add_1559_34_n_475), .B
       (count_instr[57]), .Y (inc_add_1559_34_n_470));
  AOI2BB1X1 inc_add_1559_34_g861(.A0N (count_instr[56]), .A1N
       (inc_add_1559_34_n_480), .B0 (inc_add_1559_34_n_475), .Y
       (n_6999));
  AND2X1 inc_add_1559_34_g862(.A (inc_add_1559_34_n_480), .B
       (count_instr[56]), .Y (inc_add_1559_34_n_475));
  XNOR2X1 inc_add_1559_34_g863(.A (count_instr[55]), .B
       (inc_add_1559_34_n_485), .Y (n_7000));
  NOR2BX1 inc_add_1559_34_g864(.AN (count_instr[55]), .B
       (inc_add_1559_34_n_485), .Y (inc_add_1559_34_n_480));
  OA21X1 inc_add_1559_34_g865(.A0 (count_instr[54]), .A1
       (inc_add_1559_34_n_490), .B0 (inc_add_1559_34_n_485), .Y
       (n_7001));
  NAND2X1 inc_add_1559_34_g866(.A (count_instr[54]), .B
       (inc_add_1559_34_n_490), .Y (inc_add_1559_34_n_485));
  AOI2BB1X1 inc_add_1559_34_g867(.A0N (count_instr[53]), .A1N
       (inc_add_1559_34_n_495), .B0 (inc_add_1559_34_n_490), .Y
       (n_7002));
  AND2X1 inc_add_1559_34_g868(.A (inc_add_1559_34_n_495), .B
       (count_instr[53]), .Y (inc_add_1559_34_n_490));
  XNOR2X1 inc_add_1559_34_g869(.A (count_instr[52]), .B
       (inc_add_1559_34_n_500), .Y (n_7003));
  NOR2BX1 inc_add_1559_34_g870(.AN (count_instr[52]), .B
       (inc_add_1559_34_n_500), .Y (inc_add_1559_34_n_495));
  OA21X1 inc_add_1559_34_g871(.A0 (count_instr[51]), .A1
       (inc_add_1559_34_n_505), .B0 (inc_add_1559_34_n_500), .Y
       (n_7004));
  NAND2X1 inc_add_1559_34_g872(.A (count_instr[51]), .B
       (inc_add_1559_34_n_505), .Y (inc_add_1559_34_n_500));
  AOI2BB1X1 inc_add_1559_34_g873(.A0N (count_instr[50]), .A1N
       (inc_add_1559_34_n_510), .B0 (inc_add_1559_34_n_505), .Y
       (n_7005));
  AND2X1 inc_add_1559_34_g874(.A (inc_add_1559_34_n_510), .B
       (count_instr[50]), .Y (inc_add_1559_34_n_505));
  XNOR2X1 inc_add_1559_34_g875(.A (count_instr[49]), .B
       (inc_add_1559_34_n_515), .Y (n_7006));
  NOR2BX1 inc_add_1559_34_g876(.AN (count_instr[49]), .B
       (inc_add_1559_34_n_515), .Y (inc_add_1559_34_n_510));
  OA21X1 inc_add_1559_34_g877(.A0 (count_instr[48]), .A1
       (inc_add_1559_34_n_520), .B0 (inc_add_1559_34_n_515), .Y
       (n_7007));
  NAND2X1 inc_add_1559_34_g878(.A (count_instr[48]), .B
       (inc_add_1559_34_n_520), .Y (inc_add_1559_34_n_515));
  XNOR2X1 inc_add_1559_34_g879(.A (count_instr[47]), .B
       (inc_add_1559_34_n_525), .Y (n_7008));
  NOR2BX1 inc_add_1559_34_g880(.AN (count_instr[47]), .B
       (inc_add_1559_34_n_525), .Y (inc_add_1559_34_n_520));
  OA21X1 inc_add_1559_34_g881(.A0 (count_instr[46]), .A1
       (inc_add_1559_34_n_530), .B0 (inc_add_1559_34_n_525), .Y
       (n_7009));
  NAND2X1 inc_add_1559_34_g882(.A (count_instr[46]), .B
       (inc_add_1559_34_n_530), .Y (inc_add_1559_34_n_525));
  AOI2BB1X1 inc_add_1559_34_g883(.A0N (count_instr[45]), .A1N
       (inc_add_1559_34_n_535), .B0 (inc_add_1559_34_n_530), .Y
       (n_7010));
  AND2X1 inc_add_1559_34_g884(.A (inc_add_1559_34_n_535), .B
       (count_instr[45]), .Y (inc_add_1559_34_n_530));
  XNOR2X1 inc_add_1559_34_g885(.A (count_instr[44]), .B
       (inc_add_1559_34_n_540), .Y (n_7011));
  NOR2BX1 inc_add_1559_34_g886(.AN (count_instr[44]), .B
       (inc_add_1559_34_n_540), .Y (inc_add_1559_34_n_535));
  OA21X1 inc_add_1559_34_g887(.A0 (count_instr[43]), .A1
       (inc_add_1559_34_n_545), .B0 (inc_add_1559_34_n_540), .Y
       (n_7012));
  NAND2X1 inc_add_1559_34_g888(.A (count_instr[43]), .B
       (inc_add_1559_34_n_545), .Y (inc_add_1559_34_n_540));
  AOI2BB1X1 inc_add_1559_34_g889(.A0N (count_instr[42]), .A1N
       (inc_add_1559_34_n_550), .B0 (inc_add_1559_34_n_545), .Y
       (n_7013));
  AND2X1 inc_add_1559_34_g890(.A (inc_add_1559_34_n_550), .B
       (count_instr[42]), .Y (inc_add_1559_34_n_545));
  XNOR2X1 inc_add_1559_34_g891(.A (count_instr[41]), .B
       (inc_add_1559_34_n_555), .Y (n_7014));
  NOR2BX1 inc_add_1559_34_g892(.AN (count_instr[41]), .B
       (inc_add_1559_34_n_555), .Y (inc_add_1559_34_n_550));
  XNOR2X1 inc_add_1559_34_g893(.A (count_instr[40]), .B
       (inc_add_1559_34_n_560), .Y (n_7015));
  NAND2BX1 inc_add_1559_34_g894(.AN (inc_add_1559_34_n_560), .B
       (count_instr[40]), .Y (inc_add_1559_34_n_555));
  OA21X1 inc_add_1559_34_g895(.A0 (count_instr[39]), .A1
       (inc_add_1559_34_n_565), .B0 (inc_add_1559_34_n_560), .Y
       (n_7016));
  NAND2X1 inc_add_1559_34_g896(.A (count_instr[39]), .B
       (inc_add_1559_34_n_565), .Y (inc_add_1559_34_n_560));
  AOI2BB1X1 inc_add_1559_34_g897(.A0N (count_instr[38]), .A1N
       (inc_add_1559_34_n_570), .B0 (inc_add_1559_34_n_565), .Y
       (n_7017));
  AND2X1 inc_add_1559_34_g898(.A (inc_add_1559_34_n_570), .B
       (count_instr[38]), .Y (inc_add_1559_34_n_565));
  XNOR2X1 inc_add_1559_34_g899(.A (count_instr[37]), .B
       (inc_add_1559_34_n_575), .Y (n_7018));
  NOR2BX1 inc_add_1559_34_g900(.AN (count_instr[37]), .B
       (inc_add_1559_34_n_575), .Y (inc_add_1559_34_n_570));
  OA21X1 inc_add_1559_34_g901(.A0 (count_instr[36]), .A1
       (inc_add_1559_34_n_580), .B0 (inc_add_1559_34_n_575), .Y
       (n_7019));
  NAND2X1 inc_add_1559_34_g902(.A (count_instr[36]), .B
       (inc_add_1559_34_n_580), .Y (inc_add_1559_34_n_575));
  XNOR2X1 inc_add_1559_34_g903(.A (count_instr[35]), .B
       (inc_add_1559_34_n_585), .Y (n_7020));
  NOR2BX1 inc_add_1559_34_g904(.AN (count_instr[35]), .B
       (inc_add_1559_34_n_585), .Y (inc_add_1559_34_n_580));
  OA21X1 inc_add_1559_34_g905(.A0 (count_instr[34]), .A1
       (inc_add_1559_34_n_590), .B0 (inc_add_1559_34_n_585), .Y
       (n_7021));
  NAND2X1 inc_add_1559_34_g906(.A (count_instr[34]), .B
       (inc_add_1559_34_n_590), .Y (inc_add_1559_34_n_585));
  AOI2BB1X1 inc_add_1559_34_g907(.A0N (count_instr[33]), .A1N
       (inc_add_1559_34_n_595), .B0 (inc_add_1559_34_n_590), .Y
       (n_7022));
  AND2X1 inc_add_1559_34_g908(.A (inc_add_1559_34_n_595), .B
       (count_instr[33]), .Y (inc_add_1559_34_n_590));
  XNOR2X1 inc_add_1559_34_g909(.A (count_instr[32]), .B
       (inc_add_1559_34_n_600), .Y (n_7023));
  NOR2BX1 inc_add_1559_34_g910(.AN (count_instr[32]), .B
       (inc_add_1559_34_n_600), .Y (inc_add_1559_34_n_595));
  OA21X1 inc_add_1559_34_g911(.A0 (count_instr[31]), .A1
       (inc_add_1559_34_n_605), .B0 (inc_add_1559_34_n_600), .Y
       (n_7024));
  NAND2X1 inc_add_1559_34_g912(.A (count_instr[31]), .B
       (inc_add_1559_34_n_605), .Y (inc_add_1559_34_n_600));
  AOI2BB1X1 inc_add_1559_34_g913(.A0N (count_instr[30]), .A1N
       (inc_add_1559_34_n_610), .B0 (inc_add_1559_34_n_605), .Y
       (n_7025));
  AND2X1 inc_add_1559_34_g914(.A (inc_add_1559_34_n_610), .B
       (count_instr[30]), .Y (inc_add_1559_34_n_605));
  XNOR2X1 inc_add_1559_34_g915(.A (count_instr[29]), .B
       (inc_add_1559_34_n_615), .Y (n_7026));
  NOR2BX1 inc_add_1559_34_g916(.AN (count_instr[29]), .B
       (inc_add_1559_34_n_615), .Y (inc_add_1559_34_n_610));
  OA21X1 inc_add_1559_34_g917(.A0 (count_instr[28]), .A1
       (inc_add_1559_34_n_620), .B0 (inc_add_1559_34_n_615), .Y
       (n_7027));
  NAND2X1 inc_add_1559_34_g918(.A (count_instr[28]), .B
       (inc_add_1559_34_n_620), .Y (inc_add_1559_34_n_615));
  XNOR2X1 inc_add_1559_34_g919(.A (count_instr[27]), .B
       (inc_add_1559_34_n_625), .Y (n_7028));
  NOR2BX1 inc_add_1559_34_g920(.AN (count_instr[27]), .B
       (inc_add_1559_34_n_625), .Y (inc_add_1559_34_n_620));
  OA21X1 inc_add_1559_34_g921(.A0 (count_instr[26]), .A1
       (inc_add_1559_34_n_630), .B0 (inc_add_1559_34_n_625), .Y
       (n_7029));
  NAND2X1 inc_add_1559_34_g922(.A (count_instr[26]), .B
       (inc_add_1559_34_n_630), .Y (inc_add_1559_34_n_625));
  AOI2BB1X1 inc_add_1559_34_g923(.A0N (count_instr[25]), .A1N
       (inc_add_1559_34_n_635), .B0 (inc_add_1559_34_n_630), .Y
       (n_7030));
  AND2X1 inc_add_1559_34_g924(.A (inc_add_1559_34_n_635), .B
       (count_instr[25]), .Y (inc_add_1559_34_n_630));
  AOI2BB1X1 inc_add_1559_34_g925(.A0N (count_instr[24]), .A1N
       (inc_add_1559_34_n_640), .B0 (inc_add_1559_34_n_635), .Y
       (n_7031));
  AND2X1 inc_add_1559_34_g926(.A (inc_add_1559_34_n_640), .B
       (count_instr[24]), .Y (inc_add_1559_34_n_635));
  XNOR2X1 inc_add_1559_34_g927(.A (count_instr[23]), .B
       (inc_add_1559_34_n_645), .Y (n_7032));
  NOR2BX1 inc_add_1559_34_g928(.AN (count_instr[23]), .B
       (inc_add_1559_34_n_645), .Y (inc_add_1559_34_n_640));
  OA21X1 inc_add_1559_34_g929(.A0 (count_instr[22]), .A1
       (inc_add_1559_34_n_650), .B0 (inc_add_1559_34_n_645), .Y
       (n_7033));
  NAND2X1 inc_add_1559_34_g930(.A (count_instr[22]), .B
       (inc_add_1559_34_n_650), .Y (inc_add_1559_34_n_645));
  AOI2BB1X1 inc_add_1559_34_g931(.A0N (count_instr[21]), .A1N
       (inc_add_1559_34_n_655), .B0 (inc_add_1559_34_n_650), .Y
       (n_7034));
  AND2X1 inc_add_1559_34_g932(.A (inc_add_1559_34_n_655), .B
       (count_instr[21]), .Y (inc_add_1559_34_n_650));
  XNOR2X1 inc_add_1559_34_g933(.A (count_instr[20]), .B
       (inc_add_1559_34_n_660), .Y (n_7035));
  NOR2BX1 inc_add_1559_34_g934(.AN (count_instr[20]), .B
       (inc_add_1559_34_n_660), .Y (inc_add_1559_34_n_655));
  OA21X1 inc_add_1559_34_g935(.A0 (count_instr[19]), .A1
       (inc_add_1559_34_n_665), .B0 (inc_add_1559_34_n_660), .Y
       (n_7036));
  NAND2X1 inc_add_1559_34_g936(.A (count_instr[19]), .B
       (inc_add_1559_34_n_665), .Y (inc_add_1559_34_n_660));
  AOI2BB1X1 inc_add_1559_34_g937(.A0N (count_instr[18]), .A1N
       (inc_add_1559_34_n_670), .B0 (inc_add_1559_34_n_665), .Y
       (n_7037));
  AND2X1 inc_add_1559_34_g938(.A (inc_add_1559_34_n_670), .B
       (count_instr[18]), .Y (inc_add_1559_34_n_665));
  XNOR2X1 inc_add_1559_34_g939(.A (count_instr[17]), .B
       (inc_add_1559_34_n_675), .Y (n_7038));
  NOR2BX1 inc_add_1559_34_g940(.AN (count_instr[17]), .B
       (inc_add_1559_34_n_675), .Y (inc_add_1559_34_n_670));
  XNOR2X1 inc_add_1559_34_g941(.A (count_instr[16]), .B
       (inc_add_1559_34_n_680), .Y (n_7039));
  NAND2BX1 inc_add_1559_34_g942(.AN (inc_add_1559_34_n_680), .B
       (count_instr[16]), .Y (inc_add_1559_34_n_675));
  OA21X1 inc_add_1559_34_g943(.A0 (count_instr[15]), .A1
       (inc_add_1559_34_n_685), .B0 (inc_add_1559_34_n_680), .Y
       (n_7040));
  NAND2X1 inc_add_1559_34_g944(.A (count_instr[15]), .B
       (inc_add_1559_34_n_685), .Y (inc_add_1559_34_n_680));
  AOI2BB1X1 inc_add_1559_34_g945(.A0N (count_instr[14]), .A1N
       (inc_add_1559_34_n_688), .B0 (inc_add_1559_34_n_685), .Y
       (n_7041));
  AND2X1 inc_add_1559_34_g946(.A (inc_add_1559_34_n_688), .B
       (count_instr[14]), .Y (inc_add_1559_34_n_685));
  ADDHX1 inc_add_1559_34_g947(.A (count_instr[13]), .B
       (inc_add_1559_34_n_692), .CO (inc_add_1559_34_n_688), .S
       (n_7042));
  AOI2BB1X1 inc_add_1559_34_g948(.A0N (count_instr[12]), .A1N
       (inc_add_1559_34_n_695), .B0 (inc_add_1559_34_n_692), .Y
       (n_7043));
  AND2X1 inc_add_1559_34_g949(.A (inc_add_1559_34_n_695), .B
       (count_instr[12]), .Y (inc_add_1559_34_n_692));
  ADDHX1 inc_add_1559_34_g950(.A (count_instr[11]), .B
       (inc_add_1559_34_n_699), .CO (inc_add_1559_34_n_695), .S
       (n_7044));
  AOI2BB1X1 inc_add_1559_34_g951(.A0N (count_instr[10]), .A1N
       (inc_add_1559_34_n_704), .B0 (inc_add_1559_34_n_699), .Y
       (n_7045));
  AND2X1 inc_add_1559_34_g952(.A (inc_add_1559_34_n_704), .B
       (count_instr[10]), .Y (inc_add_1559_34_n_699));
  AOI2BB1X1 inc_add_1559_34_g953(.A0N (count_instr[9]), .A1N
       (inc_add_1559_34_n_709), .B0 (inc_add_1559_34_n_704), .Y
       (n_7046));
  AND2X1 inc_add_1559_34_g954(.A (inc_add_1559_34_n_709), .B
       (count_instr[9]), .Y (inc_add_1559_34_n_704));
  XNOR2X1 inc_add_1559_34_g955(.A (count_instr[8]), .B
       (inc_add_1559_34_n_714), .Y (n_7047));
  NOR2BX1 inc_add_1559_34_g956(.AN (count_instr[8]), .B
       (inc_add_1559_34_n_714), .Y (inc_add_1559_34_n_709));
  OA21X1 inc_add_1559_34_g957(.A0 (count_instr[7]), .A1
       (inc_add_1559_34_n_719), .B0 (inc_add_1559_34_n_714), .Y
       (n_7048));
  NAND2X1 inc_add_1559_34_g958(.A (count_instr[7]), .B
       (inc_add_1559_34_n_719), .Y (inc_add_1559_34_n_714));
  AOI2BB1X1 inc_add_1559_34_g959(.A0N (count_instr[6]), .A1N
       (inc_add_1559_34_n_722), .B0 (inc_add_1559_34_n_719), .Y
       (n_7049));
  AND2X1 inc_add_1559_34_g960(.A (inc_add_1559_34_n_722), .B
       (count_instr[6]), .Y (inc_add_1559_34_n_719));
  ADDHX1 inc_add_1559_34_g961(.A (count_instr[5]), .B
       (inc_add_1559_34_n_726), .CO (inc_add_1559_34_n_722), .S
       (n_7050));
  AOI2BB1X1 inc_add_1559_34_g962(.A0N (count_instr[4]), .A1N
       (inc_add_1559_34_n_731), .B0 (inc_add_1559_34_n_726), .Y
       (n_7051));
  AND2X1 inc_add_1559_34_g963(.A (inc_add_1559_34_n_731), .B
       (count_instr[4]), .Y (inc_add_1559_34_n_726));
  AOI2BB1X1 inc_add_1559_34_g964(.A0N (count_instr[3]), .A1N
       (inc_add_1559_34_n_736), .B0 (inc_add_1559_34_n_731), .Y
       (n_7052));
  AND2X1 inc_add_1559_34_g965(.A (inc_add_1559_34_n_736), .B
       (count_instr[3]), .Y (inc_add_1559_34_n_731));
  AOI2BB1X1 inc_add_1559_34_g966(.A0N (count_instr[2]), .A1N
       (inc_add_1559_34_n_741), .B0 (inc_add_1559_34_n_736), .Y
       (n_7053));
  AND2X1 inc_add_1559_34_g967(.A (inc_add_1559_34_n_741), .B
       (count_instr[2]), .Y (inc_add_1559_34_n_736));
  AOI2BB1X1 inc_add_1559_34_g968(.A0N (count_instr[1]), .A1N
       (count_instr[0]), .B0 (inc_add_1559_34_n_741), .Y (n_7054));
  AND2X1 inc_add_1559_34_g969(.A (count_instr[0]), .B (count_instr[1]),
       .Y (inc_add_1559_34_n_741));
  XNOR2X1 inc_add_1428_40_g848(.A (count_cycle[63]), .B
       (inc_add_1428_40_n_445), .Y (n_6802));
  OA21X1 inc_add_1428_40_g849(.A0 (count_cycle[62]), .A1
       (inc_add_1428_40_n_450), .B0 (inc_add_1428_40_n_445), .Y
       (n_6801));
  NAND2X1 inc_add_1428_40_g850(.A (count_cycle[62]), .B
       (inc_add_1428_40_n_450), .Y (inc_add_1428_40_n_445));
  XNOR2X1 inc_add_1428_40_g851(.A (count_cycle[61]), .B
       (inc_add_1428_40_n_455), .Y (n_6800));
  NOR2BX1 inc_add_1428_40_g852(.AN (count_cycle[61]), .B
       (inc_add_1428_40_n_455), .Y (inc_add_1428_40_n_450));
  OA21X1 inc_add_1428_40_g853(.A0 (count_cycle[60]), .A1
       (inc_add_1428_40_n_460), .B0 (inc_add_1428_40_n_455), .Y
       (n_6799));
  NAND2X1 inc_add_1428_40_g854(.A (count_cycle[60]), .B
       (inc_add_1428_40_n_460), .Y (inc_add_1428_40_n_455));
  XNOR2X1 inc_add_1428_40_g855(.A (count_cycle[59]), .B
       (inc_add_1428_40_n_465), .Y (n_6798));
  NOR2BX1 inc_add_1428_40_g856(.AN (count_cycle[59]), .B
       (inc_add_1428_40_n_465), .Y (inc_add_1428_40_n_460));
  OA21X1 inc_add_1428_40_g857(.A0 (count_cycle[58]), .A1
       (inc_add_1428_40_n_470), .B0 (inc_add_1428_40_n_465), .Y
       (n_6797));
  NAND2X1 inc_add_1428_40_g858(.A (count_cycle[58]), .B
       (inc_add_1428_40_n_470), .Y (inc_add_1428_40_n_465));
  AOI2BB1X1 inc_add_1428_40_g859(.A0N (count_cycle[57]), .A1N
       (inc_add_1428_40_n_475), .B0 (inc_add_1428_40_n_470), .Y
       (n_6796));
  AND2X1 inc_add_1428_40_g860(.A (inc_add_1428_40_n_475), .B
       (count_cycle[57]), .Y (inc_add_1428_40_n_470));
  AOI2BB1X1 inc_add_1428_40_g861(.A0N (count_cycle[56]), .A1N
       (inc_add_1428_40_n_480), .B0 (inc_add_1428_40_n_475), .Y
       (n_6795));
  AND2X1 inc_add_1428_40_g862(.A (inc_add_1428_40_n_480), .B
       (count_cycle[56]), .Y (inc_add_1428_40_n_475));
  XNOR2X1 inc_add_1428_40_g863(.A (count_cycle[55]), .B
       (inc_add_1428_40_n_485), .Y (n_6794));
  NOR2BX1 inc_add_1428_40_g864(.AN (count_cycle[55]), .B
       (inc_add_1428_40_n_485), .Y (inc_add_1428_40_n_480));
  OA21X1 inc_add_1428_40_g865(.A0 (count_cycle[54]), .A1
       (inc_add_1428_40_n_490), .B0 (inc_add_1428_40_n_485), .Y
       (n_6793));
  NAND2X1 inc_add_1428_40_g866(.A (count_cycle[54]), .B
       (inc_add_1428_40_n_490), .Y (inc_add_1428_40_n_485));
  AOI2BB1X1 inc_add_1428_40_g867(.A0N (count_cycle[53]), .A1N
       (inc_add_1428_40_n_495), .B0 (inc_add_1428_40_n_490), .Y
       (n_6792));
  AND2X1 inc_add_1428_40_g868(.A (inc_add_1428_40_n_495), .B
       (count_cycle[53]), .Y (inc_add_1428_40_n_490));
  XNOR2X1 inc_add_1428_40_g869(.A (count_cycle[52]), .B
       (inc_add_1428_40_n_500), .Y (n_6791));
  NOR2BX1 inc_add_1428_40_g870(.AN (count_cycle[52]), .B
       (inc_add_1428_40_n_500), .Y (inc_add_1428_40_n_495));
  OA21X1 inc_add_1428_40_g871(.A0 (count_cycle[51]), .A1
       (inc_add_1428_40_n_505), .B0 (inc_add_1428_40_n_500), .Y
       (n_6790));
  NAND2X1 inc_add_1428_40_g872(.A (count_cycle[51]), .B
       (inc_add_1428_40_n_505), .Y (inc_add_1428_40_n_500));
  AOI2BB1X1 inc_add_1428_40_g873(.A0N (count_cycle[50]), .A1N
       (inc_add_1428_40_n_510), .B0 (inc_add_1428_40_n_505), .Y
       (n_6789));
  AND2X1 inc_add_1428_40_g874(.A (inc_add_1428_40_n_510), .B
       (count_cycle[50]), .Y (inc_add_1428_40_n_505));
  XNOR2X1 inc_add_1428_40_g875(.A (count_cycle[49]), .B
       (inc_add_1428_40_n_515), .Y (n_6788));
  NOR2BX1 inc_add_1428_40_g876(.AN (count_cycle[49]), .B
       (inc_add_1428_40_n_515), .Y (inc_add_1428_40_n_510));
  OA21X1 inc_add_1428_40_g877(.A0 (count_cycle[48]), .A1
       (inc_add_1428_40_n_520), .B0 (inc_add_1428_40_n_515), .Y
       (n_6787));
  NAND2X1 inc_add_1428_40_g878(.A (count_cycle[48]), .B
       (inc_add_1428_40_n_520), .Y (inc_add_1428_40_n_515));
  XNOR2X1 inc_add_1428_40_g879(.A (count_cycle[47]), .B
       (inc_add_1428_40_n_525), .Y (n_6786));
  NOR2BX1 inc_add_1428_40_g880(.AN (count_cycle[47]), .B
       (inc_add_1428_40_n_525), .Y (inc_add_1428_40_n_520));
  OA21X1 inc_add_1428_40_g881(.A0 (count_cycle[46]), .A1
       (inc_add_1428_40_n_530), .B0 (inc_add_1428_40_n_525), .Y
       (n_6785));
  NAND2X1 inc_add_1428_40_g882(.A (count_cycle[46]), .B
       (inc_add_1428_40_n_530), .Y (inc_add_1428_40_n_525));
  AOI2BB1X1 inc_add_1428_40_g883(.A0N (count_cycle[45]), .A1N
       (inc_add_1428_40_n_535), .B0 (inc_add_1428_40_n_530), .Y
       (n_6784));
  AND2X1 inc_add_1428_40_g884(.A (inc_add_1428_40_n_535), .B
       (count_cycle[45]), .Y (inc_add_1428_40_n_530));
  XNOR2X1 inc_add_1428_40_g885(.A (count_cycle[44]), .B
       (inc_add_1428_40_n_540), .Y (n_6783));
  NOR2BX1 inc_add_1428_40_g886(.AN (count_cycle[44]), .B
       (inc_add_1428_40_n_540), .Y (inc_add_1428_40_n_535));
  OA21X1 inc_add_1428_40_g887(.A0 (count_cycle[43]), .A1
       (inc_add_1428_40_n_545), .B0 (inc_add_1428_40_n_540), .Y
       (n_6782));
  NAND2X1 inc_add_1428_40_g888(.A (count_cycle[43]), .B
       (inc_add_1428_40_n_545), .Y (inc_add_1428_40_n_540));
  AOI2BB1X1 inc_add_1428_40_g889(.A0N (count_cycle[42]), .A1N
       (inc_add_1428_40_n_550), .B0 (inc_add_1428_40_n_545), .Y
       (n_6781));
  AND2X1 inc_add_1428_40_g890(.A (inc_add_1428_40_n_550), .B
       (count_cycle[42]), .Y (inc_add_1428_40_n_545));
  XNOR2X1 inc_add_1428_40_g891(.A (count_cycle[41]), .B
       (inc_add_1428_40_n_555), .Y (n_6780));
  NOR2BX1 inc_add_1428_40_g892(.AN (count_cycle[41]), .B
       (inc_add_1428_40_n_555), .Y (inc_add_1428_40_n_550));
  XNOR2X1 inc_add_1428_40_g893(.A (count_cycle[40]), .B
       (inc_add_1428_40_n_560), .Y (n_6779));
  NAND2BX1 inc_add_1428_40_g894(.AN (inc_add_1428_40_n_560), .B
       (count_cycle[40]), .Y (inc_add_1428_40_n_555));
  OA21X1 inc_add_1428_40_g895(.A0 (count_cycle[39]), .A1
       (inc_add_1428_40_n_565), .B0 (inc_add_1428_40_n_560), .Y
       (n_6778));
  NAND2X1 inc_add_1428_40_g896(.A (count_cycle[39]), .B
       (inc_add_1428_40_n_565), .Y (inc_add_1428_40_n_560));
  AOI2BB1X1 inc_add_1428_40_g897(.A0N (count_cycle[38]), .A1N
       (inc_add_1428_40_n_570), .B0 (inc_add_1428_40_n_565), .Y
       (n_6777));
  AND2X1 inc_add_1428_40_g898(.A (inc_add_1428_40_n_570), .B
       (count_cycle[38]), .Y (inc_add_1428_40_n_565));
  XNOR2X1 inc_add_1428_40_g899(.A (count_cycle[37]), .B
       (inc_add_1428_40_n_575), .Y (n_6776));
  NOR2BX1 inc_add_1428_40_g900(.AN (count_cycle[37]), .B
       (inc_add_1428_40_n_575), .Y (inc_add_1428_40_n_570));
  OA21X1 inc_add_1428_40_g901(.A0 (count_cycle[36]), .A1
       (inc_add_1428_40_n_580), .B0 (inc_add_1428_40_n_575), .Y
       (n_6775));
  NAND2X1 inc_add_1428_40_g902(.A (count_cycle[36]), .B
       (inc_add_1428_40_n_580), .Y (inc_add_1428_40_n_575));
  XNOR2X1 inc_add_1428_40_g903(.A (count_cycle[35]), .B
       (inc_add_1428_40_n_585), .Y (n_6774));
  NOR2BX1 inc_add_1428_40_g904(.AN (count_cycle[35]), .B
       (inc_add_1428_40_n_585), .Y (inc_add_1428_40_n_580));
  OA21X1 inc_add_1428_40_g905(.A0 (count_cycle[34]), .A1
       (inc_add_1428_40_n_590), .B0 (inc_add_1428_40_n_585), .Y
       (n_6773));
  NAND2X1 inc_add_1428_40_g906(.A (count_cycle[34]), .B
       (inc_add_1428_40_n_590), .Y (inc_add_1428_40_n_585));
  AOI2BB1X1 inc_add_1428_40_g907(.A0N (count_cycle[33]), .A1N
       (inc_add_1428_40_n_595), .B0 (inc_add_1428_40_n_590), .Y
       (n_6772));
  AND2X1 inc_add_1428_40_g908(.A (inc_add_1428_40_n_595), .B
       (count_cycle[33]), .Y (inc_add_1428_40_n_590));
  XNOR2X1 inc_add_1428_40_g909(.A (count_cycle[32]), .B
       (inc_add_1428_40_n_600), .Y (n_6771));
  NOR2BX1 inc_add_1428_40_g910(.AN (count_cycle[32]), .B
       (inc_add_1428_40_n_600), .Y (inc_add_1428_40_n_595));
  OA21X1 inc_add_1428_40_g911(.A0 (count_cycle[31]), .A1
       (inc_add_1428_40_n_605), .B0 (inc_add_1428_40_n_600), .Y
       (n_6770));
  NAND2X1 inc_add_1428_40_g912(.A (count_cycle[31]), .B
       (inc_add_1428_40_n_605), .Y (inc_add_1428_40_n_600));
  AOI2BB1X1 inc_add_1428_40_g913(.A0N (count_cycle[30]), .A1N
       (inc_add_1428_40_n_610), .B0 (inc_add_1428_40_n_605), .Y
       (n_6769));
  AND2X1 inc_add_1428_40_g914(.A (inc_add_1428_40_n_610), .B
       (count_cycle[30]), .Y (inc_add_1428_40_n_605));
  XNOR2X1 inc_add_1428_40_g915(.A (count_cycle[29]), .B
       (inc_add_1428_40_n_615), .Y (n_6768));
  NOR2BX1 inc_add_1428_40_g916(.AN (count_cycle[29]), .B
       (inc_add_1428_40_n_615), .Y (inc_add_1428_40_n_610));
  OA21X1 inc_add_1428_40_g917(.A0 (count_cycle[28]), .A1
       (inc_add_1428_40_n_620), .B0 (inc_add_1428_40_n_615), .Y
       (n_6767));
  NAND2X1 inc_add_1428_40_g918(.A (count_cycle[28]), .B
       (inc_add_1428_40_n_620), .Y (inc_add_1428_40_n_615));
  XNOR2X1 inc_add_1428_40_g919(.A (count_cycle[27]), .B
       (inc_add_1428_40_n_625), .Y (n_6766));
  NOR2BX1 inc_add_1428_40_g920(.AN (count_cycle[27]), .B
       (inc_add_1428_40_n_625), .Y (inc_add_1428_40_n_620));
  OA21X1 inc_add_1428_40_g921(.A0 (count_cycle[26]), .A1
       (inc_add_1428_40_n_630), .B0 (inc_add_1428_40_n_625), .Y
       (n_6765));
  NAND2X1 inc_add_1428_40_g922(.A (count_cycle[26]), .B
       (inc_add_1428_40_n_630), .Y (inc_add_1428_40_n_625));
  AOI2BB1X1 inc_add_1428_40_g923(.A0N (count_cycle[25]), .A1N
       (inc_add_1428_40_n_635), .B0 (inc_add_1428_40_n_630), .Y
       (n_6764));
  AND2X1 inc_add_1428_40_g924(.A (inc_add_1428_40_n_635), .B
       (count_cycle[25]), .Y (inc_add_1428_40_n_630));
  AOI2BB1X1 inc_add_1428_40_g925(.A0N (count_cycle[24]), .A1N
       (inc_add_1428_40_n_640), .B0 (inc_add_1428_40_n_635), .Y
       (n_6763));
  AND2X1 inc_add_1428_40_g926(.A (inc_add_1428_40_n_640), .B
       (count_cycle[24]), .Y (inc_add_1428_40_n_635));
  XNOR2X1 inc_add_1428_40_g927(.A (count_cycle[23]), .B
       (inc_add_1428_40_n_645), .Y (n_6762));
  NOR2BX1 inc_add_1428_40_g928(.AN (count_cycle[23]), .B
       (inc_add_1428_40_n_645), .Y (inc_add_1428_40_n_640));
  OA21X1 inc_add_1428_40_g929(.A0 (count_cycle[22]), .A1
       (inc_add_1428_40_n_650), .B0 (inc_add_1428_40_n_645), .Y
       (n_6761));
  NAND2X1 inc_add_1428_40_g930(.A (count_cycle[22]), .B
       (inc_add_1428_40_n_650), .Y (inc_add_1428_40_n_645));
  AOI2BB1X1 inc_add_1428_40_g931(.A0N (count_cycle[21]), .A1N
       (inc_add_1428_40_n_655), .B0 (inc_add_1428_40_n_650), .Y
       (n_6760));
  AND2X1 inc_add_1428_40_g932(.A (inc_add_1428_40_n_655), .B
       (count_cycle[21]), .Y (inc_add_1428_40_n_650));
  XNOR2X1 inc_add_1428_40_g933(.A (count_cycle[20]), .B
       (inc_add_1428_40_n_660), .Y (n_6759));
  NOR2BX1 inc_add_1428_40_g934(.AN (count_cycle[20]), .B
       (inc_add_1428_40_n_660), .Y (inc_add_1428_40_n_655));
  OA21X1 inc_add_1428_40_g935(.A0 (count_cycle[19]), .A1
       (inc_add_1428_40_n_665), .B0 (inc_add_1428_40_n_660), .Y
       (n_6758));
  NAND2X1 inc_add_1428_40_g936(.A (count_cycle[19]), .B
       (inc_add_1428_40_n_665), .Y (inc_add_1428_40_n_660));
  AOI2BB1X1 inc_add_1428_40_g937(.A0N (count_cycle[18]), .A1N
       (inc_add_1428_40_n_670), .B0 (inc_add_1428_40_n_665), .Y
       (n_6757));
  AND2X1 inc_add_1428_40_g938(.A (inc_add_1428_40_n_670), .B
       (count_cycle[18]), .Y (inc_add_1428_40_n_665));
  XNOR2X1 inc_add_1428_40_g939(.A (count_cycle[17]), .B
       (inc_add_1428_40_n_675), .Y (n_6756));
  NOR2BX1 inc_add_1428_40_g940(.AN (count_cycle[17]), .B
       (inc_add_1428_40_n_675), .Y (inc_add_1428_40_n_670));
  XNOR2X1 inc_add_1428_40_g941(.A (count_cycle[16]), .B
       (inc_add_1428_40_n_680), .Y (n_6755));
  NAND2BX1 inc_add_1428_40_g942(.AN (inc_add_1428_40_n_680), .B
       (count_cycle[16]), .Y (inc_add_1428_40_n_675));
  OA21X1 inc_add_1428_40_g943(.A0 (count_cycle[15]), .A1
       (inc_add_1428_40_n_685), .B0 (inc_add_1428_40_n_680), .Y
       (n_6754));
  NAND2X1 inc_add_1428_40_g944(.A (count_cycle[15]), .B
       (inc_add_1428_40_n_685), .Y (inc_add_1428_40_n_680));
  AOI2BB1X1 inc_add_1428_40_g945(.A0N (count_cycle[14]), .A1N
       (inc_add_1428_40_n_688), .B0 (inc_add_1428_40_n_685), .Y
       (n_6753));
  AND2X1 inc_add_1428_40_g946(.A (inc_add_1428_40_n_688), .B
       (count_cycle[14]), .Y (inc_add_1428_40_n_685));
  ADDHX1 inc_add_1428_40_g947(.A (count_cycle[13]), .B
       (inc_add_1428_40_n_692), .CO (inc_add_1428_40_n_688), .S
       (n_6752));
  AOI2BB1X1 inc_add_1428_40_g948(.A0N (count_cycle[12]), .A1N
       (inc_add_1428_40_n_695), .B0 (inc_add_1428_40_n_692), .Y
       (n_6751));
  AND2X1 inc_add_1428_40_g949(.A (inc_add_1428_40_n_695), .B
       (count_cycle[12]), .Y (inc_add_1428_40_n_692));
  ADDHX1 inc_add_1428_40_g950(.A (count_cycle[11]), .B
       (inc_add_1428_40_n_699), .CO (inc_add_1428_40_n_695), .S
       (n_6750));
  AOI2BB1X1 inc_add_1428_40_g951(.A0N (count_cycle[10]), .A1N
       (inc_add_1428_40_n_704), .B0 (inc_add_1428_40_n_699), .Y
       (n_6749));
  AND2X1 inc_add_1428_40_g952(.A (inc_add_1428_40_n_704), .B
       (count_cycle[10]), .Y (inc_add_1428_40_n_699));
  AOI2BB1X1 inc_add_1428_40_g953(.A0N (count_cycle[9]), .A1N
       (inc_add_1428_40_n_709), .B0 (inc_add_1428_40_n_704), .Y
       (n_6748));
  AND2X1 inc_add_1428_40_g954(.A (inc_add_1428_40_n_709), .B
       (count_cycle[9]), .Y (inc_add_1428_40_n_704));
  XNOR2X1 inc_add_1428_40_g955(.A (count_cycle[8]), .B
       (inc_add_1428_40_n_714), .Y (n_6747));
  NOR2BX1 inc_add_1428_40_g956(.AN (count_cycle[8]), .B
       (inc_add_1428_40_n_714), .Y (inc_add_1428_40_n_709));
  OA21X1 inc_add_1428_40_g957(.A0 (count_cycle[7]), .A1
       (inc_add_1428_40_n_719), .B0 (inc_add_1428_40_n_714), .Y
       (n_6746));
  NAND2X1 inc_add_1428_40_g958(.A (count_cycle[7]), .B
       (inc_add_1428_40_n_719), .Y (inc_add_1428_40_n_714));
  AOI2BB1X1 inc_add_1428_40_g959(.A0N (count_cycle[6]), .A1N
       (inc_add_1428_40_n_722), .B0 (inc_add_1428_40_n_719), .Y
       (n_6745));
  AND2X1 inc_add_1428_40_g960(.A (inc_add_1428_40_n_722), .B
       (count_cycle[6]), .Y (inc_add_1428_40_n_719));
  ADDHX1 inc_add_1428_40_g961(.A (count_cycle[5]), .B
       (inc_add_1428_40_n_726), .CO (inc_add_1428_40_n_722), .S
       (n_6744));
  AOI2BB1X1 inc_add_1428_40_g962(.A0N (count_cycle[4]), .A1N
       (inc_add_1428_40_n_731), .B0 (inc_add_1428_40_n_726), .Y
       (n_6743));
  AND2X1 inc_add_1428_40_g963(.A (inc_add_1428_40_n_731), .B
       (count_cycle[4]), .Y (inc_add_1428_40_n_726));
  AOI2BB1X1 inc_add_1428_40_g964(.A0N (count_cycle[3]), .A1N
       (inc_add_1428_40_n_736), .B0 (inc_add_1428_40_n_731), .Y
       (n_6742));
  AND2X1 inc_add_1428_40_g965(.A (inc_add_1428_40_n_736), .B
       (count_cycle[3]), .Y (inc_add_1428_40_n_731));
  AOI2BB1X1 inc_add_1428_40_g966(.A0N (count_cycle[2]), .A1N
       (inc_add_1428_40_n_741), .B0 (inc_add_1428_40_n_736), .Y
       (n_6741));
  AND2X1 inc_add_1428_40_g967(.A (inc_add_1428_40_n_741), .B
       (count_cycle[2]), .Y (inc_add_1428_40_n_736));
  AOI2BB1X1 inc_add_1428_40_g968(.A0N (count_cycle[1]), .A1N
       (count_cycle[0]), .B0 (inc_add_1428_40_n_741), .Y (n_6740));
  AND2X1 inc_add_1428_40_g969(.A (count_cycle[0]), .B (count_cycle[1]),
       .Y (inc_add_1428_40_n_741));
  XNOR2X1 \genblk2.pcpi_div_minus_2470_59_g500 (.A (\reg_op2[31]_9700
       ), .B (\genblk2.pcpi_div_minus_2470_59_n_324 ), .Y
       (\genblk2.pcpi_div_n_1998 ));
  AOI21X1 \genblk2.pcpi_div_minus_2470_59_g501 (.A0 (\reg_op2[30]_9699
       ), .A1 (\genblk2.pcpi_div_minus_2470_59_n_329 ), .B0
       (\genblk2.pcpi_div_minus_2470_59_n_324 ), .Y
       (\genblk2.pcpi_div_n_1999 ));
  NOR2X1 \genblk2.pcpi_div_minus_2470_59_g502 (.A (\reg_op2[30]_9699 ),
       .B (\genblk2.pcpi_div_minus_2470_59_n_329 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_324 ));
  AOI21X1 \genblk2.pcpi_div_minus_2470_59_g503 (.A0 (\reg_op2[29]_9698
       ), .A1 (\genblk2.pcpi_div_minus_2470_59_n_335 ), .B0
       (\genblk2.pcpi_div_minus_2470_59_n_330 ), .Y
       (\genblk2.pcpi_div_n_2000 ));
  INVX1 \genblk2.pcpi_div_minus_2470_59_g504 (.A
       (\genblk2.pcpi_div_minus_2470_59_n_330 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_329 ));
  NOR2X1 \genblk2.pcpi_div_minus_2470_59_g505 (.A (\reg_op2[29]_9698 ),
       .B (\genblk2.pcpi_div_minus_2470_59_n_335 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_330 ));
  OA21X1 \genblk2.pcpi_div_minus_2470_59_g506 (.A0
       (\genblk2.pcpi_div_minus_2470_59_n_479 ), .A1
       (\genblk2.pcpi_div_minus_2470_59_n_340 ), .B0
       (\genblk2.pcpi_div_minus_2470_59_n_335 ), .Y
       (\genblk2.pcpi_div_n_2001 ));
  NAND2X1 \genblk2.pcpi_div_minus_2470_59_g507 (.A
       (\genblk2.pcpi_div_minus_2470_59_n_479 ), .B
       (\genblk2.pcpi_div_minus_2470_59_n_340 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_335 ));
  AOI21X1 \genblk2.pcpi_div_minus_2470_59_g508 (.A0 (\reg_op2[27]_9696
       ), .A1 (\genblk2.pcpi_div_minus_2470_59_n_345 ), .B0
       (\genblk2.pcpi_div_minus_2470_59_n_340 ), .Y
       (\genblk2.pcpi_div_n_2002 ));
  NOR2X1 \genblk2.pcpi_div_minus_2470_59_g509 (.A (\reg_op2[27]_9696 ),
       .B (\genblk2.pcpi_div_minus_2470_59_n_345 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_340 ));
  OA21X1 \genblk2.pcpi_div_minus_2470_59_g510 (.A0
       (\genblk2.pcpi_div_minus_2470_59_n_488 ), .A1
       (\genblk2.pcpi_div_minus_2470_59_n_350 ), .B0
       (\genblk2.pcpi_div_minus_2470_59_n_345 ), .Y
       (\genblk2.pcpi_div_n_2003 ));
  NAND2X1 \genblk2.pcpi_div_minus_2470_59_g511 (.A
       (\genblk2.pcpi_div_minus_2470_59_n_488 ), .B
       (\genblk2.pcpi_div_minus_2470_59_n_350 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_345 ));
  AOI21X1 \genblk2.pcpi_div_minus_2470_59_g512 (.A0 (\reg_op2[25]_9694
       ), .A1 (\genblk2.pcpi_div_minus_2470_59_n_355 ), .B0
       (\genblk2.pcpi_div_minus_2470_59_n_350 ), .Y
       (\genblk2.pcpi_div_n_2004 ));
  NOR2X1 \genblk2.pcpi_div_minus_2470_59_g513 (.A (\reg_op2[25]_9694 ),
       .B (\genblk2.pcpi_div_minus_2470_59_n_355 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_350 ));
  OA21X1 \genblk2.pcpi_div_minus_2470_59_g514 (.A0
       (\genblk2.pcpi_div_minus_2470_59_n_483 ), .A1
       (\genblk2.pcpi_div_minus_2470_59_n_360 ), .B0
       (\genblk2.pcpi_div_minus_2470_59_n_355 ), .Y
       (\genblk2.pcpi_div_n_2005 ));
  NAND2X1 \genblk2.pcpi_div_minus_2470_59_g515 (.A
       (\genblk2.pcpi_div_minus_2470_59_n_483 ), .B
       (\genblk2.pcpi_div_minus_2470_59_n_360 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_355 ));
  AOI21X1 \genblk2.pcpi_div_minus_2470_59_g516 (.A0 (\reg_op2[23]_9692
       ), .A1 (\genblk2.pcpi_div_minus_2470_59_n_365 ), .B0
       (\genblk2.pcpi_div_minus_2470_59_n_360 ), .Y
       (\genblk2.pcpi_div_n_2006 ));
  NOR2X1 \genblk2.pcpi_div_minus_2470_59_g517 (.A (\reg_op2[23]_9692 ),
       .B (\genblk2.pcpi_div_minus_2470_59_n_365 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_360 ));
  OA21X1 \genblk2.pcpi_div_minus_2470_59_g518 (.A0
       (\genblk2.pcpi_div_minus_2470_59_n_476 ), .A1
       (\genblk2.pcpi_div_minus_2470_59_n_370 ), .B0
       (\genblk2.pcpi_div_minus_2470_59_n_365 ), .Y
       (\genblk2.pcpi_div_n_2007 ));
  NAND2X1 \genblk2.pcpi_div_minus_2470_59_g519 (.A
       (\genblk2.pcpi_div_minus_2470_59_n_476 ), .B
       (\genblk2.pcpi_div_minus_2470_59_n_370 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_365 ));
  AOI21X1 \genblk2.pcpi_div_minus_2470_59_g520 (.A0 (\reg_op2[21]_9690
       ), .A1 (\genblk2.pcpi_div_minus_2470_59_n_375 ), .B0
       (\genblk2.pcpi_div_minus_2470_59_n_370 ), .Y
       (\genblk2.pcpi_div_n_2008 ));
  NOR2X1 \genblk2.pcpi_div_minus_2470_59_g521 (.A (\reg_op2[21]_9690 ),
       .B (\genblk2.pcpi_div_minus_2470_59_n_375 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_370 ));
  OA21X1 \genblk2.pcpi_div_minus_2470_59_g522 (.A0
       (\genblk2.pcpi_div_minus_2470_59_n_500 ), .A1
       (\genblk2.pcpi_div_minus_2470_59_n_380 ), .B0
       (\genblk2.pcpi_div_minus_2470_59_n_375 ), .Y
       (\genblk2.pcpi_div_n_2009 ));
  NAND2X1 \genblk2.pcpi_div_minus_2470_59_g523 (.A
       (\genblk2.pcpi_div_minus_2470_59_n_500 ), .B
       (\genblk2.pcpi_div_minus_2470_59_n_380 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_375 ));
  AOI21X1 \genblk2.pcpi_div_minus_2470_59_g524 (.A0 (\reg_op2[19]_9688
       ), .A1 (\genblk2.pcpi_div_minus_2470_59_n_385 ), .B0
       (\genblk2.pcpi_div_minus_2470_59_n_380 ), .Y
       (\genblk2.pcpi_div_n_2010 ));
  NOR2X1 \genblk2.pcpi_div_minus_2470_59_g525 (.A (\reg_op2[19]_9688 ),
       .B (\genblk2.pcpi_div_minus_2470_59_n_385 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_380 ));
  OA21X1 \genblk2.pcpi_div_minus_2470_59_g526 (.A0
       (\genblk2.pcpi_div_minus_2470_59_n_485 ), .A1
       (\genblk2.pcpi_div_minus_2470_59_n_390 ), .B0
       (\genblk2.pcpi_div_minus_2470_59_n_385 ), .Y
       (\genblk2.pcpi_div_n_2011 ));
  NAND2X1 \genblk2.pcpi_div_minus_2470_59_g527 (.A
       (\genblk2.pcpi_div_minus_2470_59_n_485 ), .B
       (\genblk2.pcpi_div_minus_2470_59_n_390 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_385 ));
  AOI21X1 \genblk2.pcpi_div_minus_2470_59_g528 (.A0 (\reg_op2[17]_9686
       ), .A1 (\genblk2.pcpi_div_minus_2470_59_n_395 ), .B0
       (\genblk2.pcpi_div_minus_2470_59_n_390 ), .Y
       (\genblk2.pcpi_div_n_2012 ));
  NOR2X1 \genblk2.pcpi_div_minus_2470_59_g529 (.A (\reg_op2[17]_9686 ),
       .B (\genblk2.pcpi_div_minus_2470_59_n_395 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_390 ));
  OA21X1 \genblk2.pcpi_div_minus_2470_59_g530 (.A0
       (\genblk2.pcpi_div_minus_2470_59_n_481 ), .A1
       (\genblk2.pcpi_div_minus_2470_59_n_400 ), .B0
       (\genblk2.pcpi_div_minus_2470_59_n_395 ), .Y
       (\genblk2.pcpi_div_n_2013 ));
  NAND2X1 \genblk2.pcpi_div_minus_2470_59_g531 (.A
       (\genblk2.pcpi_div_minus_2470_59_n_481 ), .B
       (\genblk2.pcpi_div_minus_2470_59_n_400 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_395 ));
  AOI21X1 \genblk2.pcpi_div_minus_2470_59_g532 (.A0 (\reg_op2[15]_9684
       ), .A1 (\genblk2.pcpi_div_minus_2470_59_n_405 ), .B0
       (\genblk2.pcpi_div_minus_2470_59_n_400 ), .Y
       (\genblk2.pcpi_div_n_2014 ));
  NOR2X1 \genblk2.pcpi_div_minus_2470_59_g533 (.A (\reg_op2[15]_9684 ),
       .B (\genblk2.pcpi_div_minus_2470_59_n_405 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_400 ));
  OA21X1 \genblk2.pcpi_div_minus_2470_59_g534 (.A0
       (\genblk2.pcpi_div_minus_2470_59_n_499 ), .A1
       (\genblk2.pcpi_div_minus_2470_59_n_410 ), .B0
       (\genblk2.pcpi_div_minus_2470_59_n_405 ), .Y
       (\genblk2.pcpi_div_n_2015 ));
  NAND2X1 \genblk2.pcpi_div_minus_2470_59_g535 (.A
       (\genblk2.pcpi_div_minus_2470_59_n_499 ), .B
       (\genblk2.pcpi_div_minus_2470_59_n_410 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_405 ));
  AOI21X1 \genblk2.pcpi_div_minus_2470_59_g536 (.A0 (\reg_op2[13]_9682
       ), .A1 (\genblk2.pcpi_div_minus_2470_59_n_415 ), .B0
       (\genblk2.pcpi_div_minus_2470_59_n_410 ), .Y
       (\genblk2.pcpi_div_n_2016 ));
  NOR2X1 \genblk2.pcpi_div_minus_2470_59_g537 (.A (\reg_op2[13]_9682 ),
       .B (\genblk2.pcpi_div_minus_2470_59_n_415 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_410 ));
  OA21X1 \genblk2.pcpi_div_minus_2470_59_g538 (.A0
       (\genblk2.pcpi_div_minus_2470_59_n_498 ), .A1
       (\genblk2.pcpi_div_minus_2470_59_n_420 ), .B0
       (\genblk2.pcpi_div_minus_2470_59_n_415 ), .Y
       (\genblk2.pcpi_div_n_2017 ));
  NAND2X1 \genblk2.pcpi_div_minus_2470_59_g539 (.A
       (\genblk2.pcpi_div_minus_2470_59_n_498 ), .B
       (\genblk2.pcpi_div_minus_2470_59_n_420 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_415 ));
  AOI21X1 \genblk2.pcpi_div_minus_2470_59_g540 (.A0 (\reg_op2[11]_9680
       ), .A1 (\genblk2.pcpi_div_minus_2470_59_n_425 ), .B0
       (\genblk2.pcpi_div_minus_2470_59_n_420 ), .Y
       (\genblk2.pcpi_div_n_2018 ));
  NOR2X1 \genblk2.pcpi_div_minus_2470_59_g541 (.A (\reg_op2[11]_9680 ),
       .B (\genblk2.pcpi_div_minus_2470_59_n_425 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_420 ));
  OA21X1 \genblk2.pcpi_div_minus_2470_59_g542 (.A0
       (\genblk2.pcpi_div_minus_2470_59_n_502 ), .A1
       (\genblk2.pcpi_div_minus_2470_59_n_430 ), .B0
       (\genblk2.pcpi_div_minus_2470_59_n_425 ), .Y
       (\genblk2.pcpi_div_n_2019 ));
  NAND2X1 \genblk2.pcpi_div_minus_2470_59_g543 (.A
       (\genblk2.pcpi_div_minus_2470_59_n_502 ), .B
       (\genblk2.pcpi_div_minus_2470_59_n_430 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_425 ));
  AOI21X1 \genblk2.pcpi_div_minus_2470_59_g544 (.A0 (\reg_op2[9]_9678
       ), .A1 (\genblk2.pcpi_div_minus_2470_59_n_435 ), .B0
       (\genblk2.pcpi_div_minus_2470_59_n_430 ), .Y
       (\genblk2.pcpi_div_n_2020 ));
  NOR2X1 \genblk2.pcpi_div_minus_2470_59_g545 (.A (\reg_op2[9]_9678 ),
       .B (\genblk2.pcpi_div_minus_2470_59_n_435 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_430 ));
  OA21X1 \genblk2.pcpi_div_minus_2470_59_g546 (.A0
       (\genblk2.pcpi_div_minus_2470_59_n_492 ), .A1
       (\genblk2.pcpi_div_minus_2470_59_n_440 ), .B0
       (\genblk2.pcpi_div_minus_2470_59_n_435 ), .Y
       (\genblk2.pcpi_div_n_2021 ));
  NAND2X1 \genblk2.pcpi_div_minus_2470_59_g547 (.A
       (\genblk2.pcpi_div_minus_2470_59_n_492 ), .B
       (\genblk2.pcpi_div_minus_2470_59_n_440 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_435 ));
  AOI21X1 \genblk2.pcpi_div_minus_2470_59_g548 (.A0 (\reg_op2[7]_9676
       ), .A1 (\genblk2.pcpi_div_minus_2470_59_n_445 ), .B0
       (\genblk2.pcpi_div_minus_2470_59_n_440 ), .Y
       (\genblk2.pcpi_div_n_2022 ));
  NOR2X1 \genblk2.pcpi_div_minus_2470_59_g549 (.A (\reg_op2[7]_9676 ),
       .B (\genblk2.pcpi_div_minus_2470_59_n_445 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_440 ));
  OA21X1 \genblk2.pcpi_div_minus_2470_59_g550 (.A0
       (\genblk2.pcpi_div_minus_2470_59_n_474 ), .A1
       (\genblk2.pcpi_div_minus_2470_59_n_450 ), .B0
       (\genblk2.pcpi_div_minus_2470_59_n_445 ), .Y
       (\genblk2.pcpi_div_n_2023 ));
  NAND2X1 \genblk2.pcpi_div_minus_2470_59_g551 (.A
       (\genblk2.pcpi_div_minus_2470_59_n_474 ), .B
       (\genblk2.pcpi_div_minus_2470_59_n_450 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_445 ));
  AOI21X1 \genblk2.pcpi_div_minus_2470_59_g552 (.A0 (\reg_op2[5]_9674
       ), .A1 (\genblk2.pcpi_div_minus_2470_59_n_455 ), .B0
       (\genblk2.pcpi_div_minus_2470_59_n_450 ), .Y
       (\genblk2.pcpi_div_n_2024 ));
  NOR2X1 \genblk2.pcpi_div_minus_2470_59_g553 (.A (\reg_op2[5]_9674 ),
       .B (\genblk2.pcpi_div_minus_2470_59_n_455 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_450 ));
  OA21X1 \genblk2.pcpi_div_minus_2470_59_g554 (.A0
       (\genblk2.pcpi_div_minus_2470_59_n_477 ), .A1
       (\genblk2.pcpi_div_minus_2470_59_n_460 ), .B0
       (\genblk2.pcpi_div_minus_2470_59_n_455 ), .Y
       (\genblk2.pcpi_div_n_2025 ));
  NAND2X1 \genblk2.pcpi_div_minus_2470_59_g555 (.A
       (\genblk2.pcpi_div_minus_2470_59_n_477 ), .B
       (\genblk2.pcpi_div_minus_2470_59_n_460 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_455 ));
  AOI21X1 \genblk2.pcpi_div_minus_2470_59_g556 (.A0 (\reg_op2[3]_9672
       ), .A1 (\genblk2.pcpi_div_minus_2470_59_n_465 ), .B0
       (\genblk2.pcpi_div_minus_2470_59_n_460 ), .Y
       (\genblk2.pcpi_div_n_2026 ));
  NOR2X1 \genblk2.pcpi_div_minus_2470_59_g557 (.A (\reg_op2[3]_9672 ),
       .B (\genblk2.pcpi_div_minus_2470_59_n_465 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_460 ));
  OA21X1 \genblk2.pcpi_div_minus_2470_59_g558 (.A0
       (\genblk2.pcpi_div_minus_2470_59_n_487 ), .A1
       (\genblk2.pcpi_div_minus_2470_59_n_470 ), .B0
       (\genblk2.pcpi_div_minus_2470_59_n_465 ), .Y
       (\genblk2.pcpi_div_n_2027 ));
  NAND2X1 \genblk2.pcpi_div_minus_2470_59_g559 (.A
       (\genblk2.pcpi_div_minus_2470_59_n_487 ), .B
       (\genblk2.pcpi_div_minus_2470_59_n_470 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_465 ));
  AOI21X1 \genblk2.pcpi_div_minus_2470_59_g560 (.A0 (\reg_op2[1]_9670
       ), .A1 (\reg_op2[0]_9669 ), .B0
       (\genblk2.pcpi_div_minus_2470_59_n_470 ), .Y
       (\genblk2.pcpi_div_n_2028 ));
  NOR2X1 \genblk2.pcpi_div_minus_2470_59_g561 (.A (\reg_op2[1]_9670 ),
       .B (\reg_op2[0]_9669 ), .Y
       (\genblk2.pcpi_div_minus_2470_59_n_470 ));
  INVX1 \genblk2.pcpi_div_minus_2470_59_g563 (.A (\reg_op2[22]_9691 ),
       .Y (\genblk2.pcpi_div_minus_2470_59_n_476 ));
  XNOR2X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g500 (.A
       (\genblk2.pcpi_div_n_2110 ), .B
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_323 ), .Y
       (\genblk2.pcpi_div_n_2142 ));
  AOI21X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g501 (.A0
       (\genblk2.pcpi_div_n_2111 ), .A1
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_328 ), .B0
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_323 ), .Y
       (\genblk2.pcpi_div_n_2143 ));
  NOR2X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g502 (.A
       (\genblk2.pcpi_div_n_2111 ), .B
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_328 ), .Y
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_323 ));
  AOI21X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g503 (.A0
       (\genblk2.pcpi_div_n_2112 ), .A1
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_334 ), .B0
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_329 ), .Y
       (\genblk2.pcpi_div_n_2144 ));
  INVX1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g504 (.A
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_329 ), .Y
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_328 ));
  NOR2X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g505 (.A
       (\genblk2.pcpi_div_n_2112 ), .B
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_334 ), .Y
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_329 ));
  OA21X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g506 (.A0
       (n_11698), .A1
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_339 ), .B0
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_334 ), .Y
       (\genblk2.pcpi_div_n_2145 ));
  NAND2X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g507 (.A
       (n_11698), .B
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_339 ), .Y
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_334 ));
  AOI21X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g508 (.A0
       (\genblk2.pcpi_div_n_2114 ), .A1
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_344 ), .B0
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_339 ), .Y
       (\genblk2.pcpi_div_n_2146 ));
  NOR2X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g509 (.A
       (\genblk2.pcpi_div_n_2114 ), .B
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_344 ), .Y
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_339 ));
  OA21X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g510 (.A0
       (n_11702), .A1
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_349 ), .B0
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_344 ), .Y
       (\genblk2.pcpi_div_n_2147 ));
  NAND2X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g511 (.A
       (n_11702), .B
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_349 ), .Y
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_344 ));
  AOI21X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g512 (.A0
       (\genblk2.pcpi_div_n_2116 ), .A1
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_354 ), .B0
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_349 ), .Y
       (\genblk2.pcpi_div_n_2148 ));
  NOR2X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g513 (.A
       (\genblk2.pcpi_div_n_2116 ), .B
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_354 ), .Y
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_349 ));
  OA21X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g514 (.A0
       (n_11705), .A1
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_359 ), .B0
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_354 ), .Y
       (\genblk2.pcpi_div_n_2149 ));
  NAND2X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g515 (.A
       (n_11705), .B
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_359 ), .Y
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_354 ));
  AOI21X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g516 (.A0
       (\genblk2.pcpi_div_n_2118 ), .A1
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_364 ), .B0
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_359 ), .Y
       (\genblk2.pcpi_div_n_2150 ));
  NOR2X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g517 (.A
       (\genblk2.pcpi_div_n_2118 ), .B
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_364 ), .Y
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_359 ));
  OA21X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g518 (.A0
       (n_11699), .A1
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_369 ), .B0
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_364 ), .Y
       (\genblk2.pcpi_div_n_2151 ));
  NAND2X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g519 (.A
       (n_11699), .B
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_369 ), .Y
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_364 ));
  AOI21X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g520 (.A0
       (\genblk2.pcpi_div_n_2120 ), .A1
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_374 ), .B0
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_369 ), .Y
       (\genblk2.pcpi_div_n_2152 ));
  NOR2X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g521 (.A
       (\genblk2.pcpi_div_n_2120 ), .B
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_374 ), .Y
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_369 ));
  OA21X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g522 (.A0
       (n_11703), .A1
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_379 ), .B0
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_374 ), .Y
       (\genblk2.pcpi_div_n_2153 ));
  NAND2X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g523 (.A
       (n_11703), .B
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_379 ), .Y
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_374 ));
  AOI21X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g524 (.A0
       (\genblk2.pcpi_div_n_2122 ), .A1
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_384 ), .B0
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_379 ), .Y
       (\genblk2.pcpi_div_n_2154 ));
  NOR2X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g525 (.A
       (\genblk2.pcpi_div_n_2122 ), .B
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_384 ), .Y
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_379 ));
  OA21X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g526 (.A0
       (n_11697), .A1
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_389 ), .B0
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_384 ), .Y
       (\genblk2.pcpi_div_n_2155 ));
  NAND2X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g527 (.A
       (n_11697), .B
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_389 ), .Y
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_384 ));
  AOI21X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g528 (.A0
       (\genblk2.pcpi_div_n_2124 ), .A1
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_394 ), .B0
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_389 ), .Y
       (\genblk2.pcpi_div_n_2156 ));
  NOR2X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g529 (.A
       (\genblk2.pcpi_div_n_2124 ), .B
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_394 ), .Y
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_389 ));
  OA21X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g530 (.A0
       (n_11696), .A1
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_399 ), .B0
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_394 ), .Y
       (\genblk2.pcpi_div_n_2157 ));
  NAND2X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g531 (.A
       (n_11696), .B
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_399 ), .Y
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_394 ));
  AOI21X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g532 (.A0
       (\genblk2.pcpi_div_n_2126 ), .A1
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_404 ), .B0
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_399 ), .Y
       (\genblk2.pcpi_div_n_2158 ));
  NOR2X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g533 (.A
       (\genblk2.pcpi_div_n_2126 ), .B
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_404 ), .Y
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_399 ));
  OA21X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g534 (.A0
       (n_11692), .A1
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_409 ), .B0
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_404 ), .Y
       (\genblk2.pcpi_div_n_2159 ));
  NAND2X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g535 (.A
       (n_11692), .B
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_409 ), .Y
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_404 ));
  AOI21X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g536 (.A0
       (\genblk2.pcpi_div_n_2128 ), .A1
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_414 ), .B0
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_409 ), .Y
       (\genblk2.pcpi_div_n_2160 ));
  NOR2X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g537 (.A
       (\genblk2.pcpi_div_n_2128 ), .B
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_414 ), .Y
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_409 ));
  OA21X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g538 (.A0
       (n_11704), .A1
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_419 ), .B0
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_414 ), .Y
       (\genblk2.pcpi_div_n_2161 ));
  NAND2X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g539 (.A
       (n_11704), .B
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_419 ), .Y
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_414 ));
  AOI21X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g540 (.A0
       (\genblk2.pcpi_div_n_2130 ), .A1
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_424 ), .B0
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_419 ), .Y
       (\genblk2.pcpi_div_n_2162 ));
  NOR2X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g541 (.A
       (\genblk2.pcpi_div_n_2130 ), .B
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_424 ), .Y
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_419 ));
  OA21X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g542 (.A0
       (n_11693), .A1
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_429 ), .B0
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_424 ), .Y
       (\genblk2.pcpi_div_n_2163 ));
  NAND2X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g543 (.A
       (n_11693), .B
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_429 ), .Y
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_424 ));
  AOI21X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g544 (.A0
       (\genblk2.pcpi_div_n_2132 ), .A1
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_434 ), .B0
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_429 ), .Y
       (\genblk2.pcpi_div_n_2164 ));
  NOR2X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g545 (.A
       (\genblk2.pcpi_div_n_2132 ), .B
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_434 ), .Y
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_429 ));
  OA21X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g546 (.A0
       (n_11695), .A1
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_439 ), .B0
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_434 ), .Y
       (\genblk2.pcpi_div_n_2165 ));
  NAND2X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g547 (.A
       (n_11695), .B
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_439 ), .Y
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_434 ));
  AOI21X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g548 (.A0
       (\genblk2.pcpi_div_n_2134 ), .A1
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_444 ), .B0
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_439 ), .Y
       (\genblk2.pcpi_div_n_2166 ));
  NOR2X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g549 (.A
       (\genblk2.pcpi_div_n_2134 ), .B
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_444 ), .Y
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_439 ));
  OA21X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g550 (.A0
       (n_11694), .A1
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_449 ), .B0
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_444 ), .Y
       (\genblk2.pcpi_div_n_2167 ));
  NAND2X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g551 (.A
       (n_11694), .B
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_449 ), .Y
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_444 ));
  AOI21X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g552 (.A0
       (\genblk2.pcpi_div_n_2136 ), .A1
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_454 ), .B0
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_449 ), .Y
       (\genblk2.pcpi_div_n_2168 ));
  NOR2X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g553 (.A
       (\genblk2.pcpi_div_n_2136 ), .B
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_454 ), .Y
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_449 ));
  OA21X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g554 (.A0
       (n_11701), .A1
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_459 ), .B0
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_454 ), .Y
       (\genblk2.pcpi_div_n_2169 ));
  NAND2X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g555 (.A
       (n_11701), .B
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_459 ), .Y
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_454 ));
  AOI21X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g556 (.A0
       (\genblk2.pcpi_div_n_2138 ), .A1
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_464 ), .B0
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_459 ), .Y
       (\genblk2.pcpi_div_n_2170 ));
  NOR2X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g557 (.A
       (\genblk2.pcpi_div_n_2138 ), .B
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_464 ), .Y
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_459 ));
  OA21X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g558 (.A0
       (n_11700), .A1
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_469 ), .B0
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_464 ), .Y
       (\genblk2.pcpi_div_n_2171 ));
  NAND2X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g559 (.A
       (n_11700), .B
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_469 ), .Y
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_464 ));
  AOI21X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g560 (.A0
       (\genblk2.pcpi_div_n_2140 ), .A1 (\genblk2.pcpi_div_n_578 ), .B0
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_469 ), .Y
       (\genblk2.pcpi_div_n_2172 ));
  NOR2X1 \genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_g561 (.A
       (\genblk2.pcpi_div_n_2140 ), .B (\genblk2.pcpi_div_n_578 ), .Y
       (\genblk2.pcpi_div_minus_2490_26_Y_minus_2488_26_n_469 ));
  XNOR2X1 sub_1235_38_Y_add_1235_58_g2863(.A
       (sub_1235_38_Y_add_1235_58_n_1407), .B
       (sub_1235_38_Y_add_1235_58_n_1346), .Y (n_6656));
  ADDFX1 sub_1235_38_Y_add_1235_58_g2864(.A (\reg_op1[30]_9667 ), .B
       (sub_1235_38_Y_add_1235_58_n_1437), .CI
       (sub_1235_38_Y_add_1235_58_n_1348), .CO
       (sub_1235_38_Y_add_1235_58_n_1346), .S (n_6655));
  ADDFX1 sub_1235_38_Y_add_1235_58_g2865(.A (\reg_op1[29]_9666 ), .B
       (sub_1235_38_Y_add_1235_58_n_1431), .CI
       (sub_1235_38_Y_add_1235_58_n_1350), .CO
       (sub_1235_38_Y_add_1235_58_n_1348), .S (n_6654));
  ADDFX1 sub_1235_38_Y_add_1235_58_g2866(.A (\reg_op1[28]_9665 ), .B
       (sub_1235_38_Y_add_1235_58_n_1410), .CI
       (sub_1235_38_Y_add_1235_58_n_1352), .CO
       (sub_1235_38_Y_add_1235_58_n_1350), .S (n_6653));
  ADDFX1 sub_1235_38_Y_add_1235_58_g2867(.A (\reg_op1[27]_9664 ), .B
       (sub_1235_38_Y_add_1235_58_n_1412), .CI
       (sub_1235_38_Y_add_1235_58_n_1354), .CO
       (sub_1235_38_Y_add_1235_58_n_1352), .S (n_6652));
  ADDFX1 sub_1235_38_Y_add_1235_58_g2868(.A (\reg_op1[26]_9663 ), .B
       (sub_1235_38_Y_add_1235_58_n_1423), .CI
       (sub_1235_38_Y_add_1235_58_n_1356), .CO
       (sub_1235_38_Y_add_1235_58_n_1354), .S (n_6651));
  ADDFX1 sub_1235_38_Y_add_1235_58_g2869(.A (\reg_op1[25]_9662 ), .B
       (sub_1235_38_Y_add_1235_58_n_1439), .CI
       (sub_1235_38_Y_add_1235_58_n_1358), .CO
       (sub_1235_38_Y_add_1235_58_n_1356), .S (n_6650));
  ADDFX1 sub_1235_38_Y_add_1235_58_g2870(.A (\reg_op1[24]_9661 ), .B
       (sub_1235_38_Y_add_1235_58_n_1416), .CI
       (sub_1235_38_Y_add_1235_58_n_1360), .CO
       (sub_1235_38_Y_add_1235_58_n_1358), .S (n_6649));
  ADDFX1 sub_1235_38_Y_add_1235_58_g2871(.A (\reg_op1[23]_9660 ), .B
       (sub_1235_38_Y_add_1235_58_n_1434), .CI
       (sub_1235_38_Y_add_1235_58_n_1362), .CO
       (sub_1235_38_Y_add_1235_58_n_1360), .S (n_6648));
  ADDFX1 sub_1235_38_Y_add_1235_58_g2872(.A (\reg_op1[22]_9659 ), .B
       (sub_1235_38_Y_add_1235_58_n_1427), .CI
       (sub_1235_38_Y_add_1235_58_n_1364), .CO
       (sub_1235_38_Y_add_1235_58_n_1362), .S (n_6647));
  ADDFX1 sub_1235_38_Y_add_1235_58_g2873(.A (\reg_op1[21]_9658 ), .B
       (sub_1235_38_Y_add_1235_58_n_1421), .CI
       (sub_1235_38_Y_add_1235_58_n_1366), .CO
       (sub_1235_38_Y_add_1235_58_n_1364), .S (n_6646));
  ADDFX1 sub_1235_38_Y_add_1235_58_g2874(.A (\reg_op1[20]_9657 ), .B
       (sub_1235_38_Y_add_1235_58_n_1420), .CI
       (sub_1235_38_Y_add_1235_58_n_1368), .CO
       (sub_1235_38_Y_add_1235_58_n_1366), .S (n_6645));
  ADDFX1 sub_1235_38_Y_add_1235_58_g2875(.A (\reg_op1[19]_9656 ), .B
       (sub_1235_38_Y_add_1235_58_n_1414), .CI
       (sub_1235_38_Y_add_1235_58_n_1370), .CO
       (sub_1235_38_Y_add_1235_58_n_1368), .S (n_6644));
  ADDFX1 sub_1235_38_Y_add_1235_58_g2876(.A (\reg_op1[18]_9655 ), .B
       (sub_1235_38_Y_add_1235_58_n_1440), .CI
       (sub_1235_38_Y_add_1235_58_n_1372), .CO
       (sub_1235_38_Y_add_1235_58_n_1370), .S (n_6643));
  ADDFX1 sub_1235_38_Y_add_1235_58_g2877(.A (\reg_op1[17]_9654 ), .B
       (sub_1235_38_Y_add_1235_58_n_1433), .CI
       (sub_1235_38_Y_add_1235_58_n_1374), .CO
       (sub_1235_38_Y_add_1235_58_n_1372), .S (n_6642));
  ADDFX1 sub_1235_38_Y_add_1235_58_g2878(.A (\reg_op1[16]_9653 ), .B
       (sub_1235_38_Y_add_1235_58_n_1418), .CI
       (sub_1235_38_Y_add_1235_58_n_1376), .CO
       (sub_1235_38_Y_add_1235_58_n_1374), .S (n_6641));
  ADDFX1 sub_1235_38_Y_add_1235_58_g2879(.A (\reg_op1[15]_9652 ), .B
       (sub_1235_38_Y_add_1235_58_n_1432), .CI
       (sub_1235_38_Y_add_1235_58_n_1378), .CO
       (sub_1235_38_Y_add_1235_58_n_1376), .S (n_6640));
  ADDFX1 sub_1235_38_Y_add_1235_58_g2880(.A (\reg_op1[14]_9651 ), .B
       (sub_1235_38_Y_add_1235_58_n_1424), .CI
       (sub_1235_38_Y_add_1235_58_n_1380), .CO
       (sub_1235_38_Y_add_1235_58_n_1378), .S (n_6639));
  ADDFX1 sub_1235_38_Y_add_1235_58_g2881(.A (\reg_op1[13]_9650 ), .B
       (sub_1235_38_Y_add_1235_58_n_1441), .CI
       (sub_1235_38_Y_add_1235_58_n_1382), .CO
       (sub_1235_38_Y_add_1235_58_n_1380), .S (n_6638));
  ADDFX1 sub_1235_38_Y_add_1235_58_g2882(.A (\reg_op1[12]_9649 ), .B
       (sub_1235_38_Y_add_1235_58_n_1428), .CI
       (sub_1235_38_Y_add_1235_58_n_1384), .CO
       (sub_1235_38_Y_add_1235_58_n_1382), .S (n_6637));
  ADDFX1 sub_1235_38_Y_add_1235_58_g2883(.A (\reg_op1[11]_9648 ), .B
       (sub_1235_38_Y_add_1235_58_n_1429), .CI
       (sub_1235_38_Y_add_1235_58_n_1386), .CO
       (sub_1235_38_Y_add_1235_58_n_1384), .S (n_6636));
  ADDFX1 sub_1235_38_Y_add_1235_58_g2884(.A (\reg_op1[10]_9647 ), .B
       (sub_1235_38_Y_add_1235_58_n_1408), .CI
       (sub_1235_38_Y_add_1235_58_n_1388), .CO
       (sub_1235_38_Y_add_1235_58_n_1386), .S (n_6635));
  ADDFX1 sub_1235_38_Y_add_1235_58_g2885(.A (\reg_op1[9]_9646 ), .B
       (sub_1235_38_Y_add_1235_58_n_1419), .CI
       (sub_1235_38_Y_add_1235_58_n_1390), .CO
       (sub_1235_38_Y_add_1235_58_n_1388), .S (n_6634));
  ADDFX1 sub_1235_38_Y_add_1235_58_g2886(.A (\reg_op1[8]_9645 ), .B
       (sub_1235_38_Y_add_1235_58_n_1435), .CI
       (sub_1235_38_Y_add_1235_58_n_1392), .CO
       (sub_1235_38_Y_add_1235_58_n_1390), .S (n_6633));
  ADDFX1 sub_1235_38_Y_add_1235_58_g2887(.A (\reg_op1[7]_9644 ), .B
       (sub_1235_38_Y_add_1235_58_n_1415), .CI
       (sub_1235_38_Y_add_1235_58_n_1394), .CO
       (sub_1235_38_Y_add_1235_58_n_1392), .S (n_6632));
  ADDFX1 sub_1235_38_Y_add_1235_58_g2888(.A (\reg_op1[6]_9643 ), .B
       (sub_1235_38_Y_add_1235_58_n_1436), .CI
       (sub_1235_38_Y_add_1235_58_n_1396), .CO
       (sub_1235_38_Y_add_1235_58_n_1394), .S (n_6631));
  ADDFX1 sub_1235_38_Y_add_1235_58_g2889(.A (\reg_op1[5]_9642 ), .B
       (sub_1235_38_Y_add_1235_58_n_1438), .CI
       (sub_1235_38_Y_add_1235_58_n_1398), .CO
       (sub_1235_38_Y_add_1235_58_n_1396), .S (n_6630));
  ADDFX1 sub_1235_38_Y_add_1235_58_g2890(.A (\reg_op1[4]_9641 ), .B
       (sub_1235_38_Y_add_1235_58_n_1426), .CI
       (sub_1235_38_Y_add_1235_58_n_1400), .CO
       (sub_1235_38_Y_add_1235_58_n_1398), .S (n_6629));
  ADDFX1 sub_1235_38_Y_add_1235_58_g2891(.A (\reg_op1[3]_9640 ), .B
       (sub_1235_38_Y_add_1235_58_n_1422), .CI
       (sub_1235_38_Y_add_1235_58_n_1402), .CO
       (sub_1235_38_Y_add_1235_58_n_1400), .S (n_6628));
  ADDFX1 sub_1235_38_Y_add_1235_58_g2892(.A (\reg_op1[2]_9639 ), .B
       (sub_1235_38_Y_add_1235_58_n_1413), .CI
       (sub_1235_38_Y_add_1235_58_n_1404), .CO
       (sub_1235_38_Y_add_1235_58_n_1402), .S (n_6627));
  ADDFX1 sub_1235_38_Y_add_1235_58_g2893(.A (\reg_op1[1]_9638 ), .B
       (sub_1235_38_Y_add_1235_58_n_1417), .CI
       (sub_1235_38_Y_add_1235_58_n_1406), .CO
       (sub_1235_38_Y_add_1235_58_n_1404), .S (n_6626));
  ADDFX1 sub_1235_38_Y_add_1235_58_g2894(.A (reg_op1[0]), .B
       (instr_sub), .CI (sub_1235_38_Y_add_1235_58_n_1425), .CO
       (sub_1235_38_Y_add_1235_58_n_1406), .S (n_6625));
  XNOR2X1 sub_1235_38_Y_add_1235_58_g2895(.A (\reg_op1[31]_9668 ), .B
       (sub_1235_38_Y_add_1235_58_n_1430), .Y
       (sub_1235_38_Y_add_1235_58_n_1407));
  MX2X1 sub_1235_38_Y_add_1235_58_g2896(.A (instr_sub), .B
       (sub_1235_38_Y_add_1235_58_n_1443), .S0 (\reg_op2[10]_9679 ), .Y
       (sub_1235_38_Y_add_1235_58_n_1408));
  MX2X1 sub_1235_38_Y_add_1235_58_g2897(.A (instr_sub), .B
       (sub_1235_38_Y_add_1235_58_n_1443), .S0 (\reg_op2[28]_9697 ), .Y
       (sub_1235_38_Y_add_1235_58_n_1410));
  MX2X1 sub_1235_38_Y_add_1235_58_g2898(.A (instr_sub), .B
       (sub_1235_38_Y_add_1235_58_n_1443), .S0 (\reg_op2[27]_9696 ), .Y
       (sub_1235_38_Y_add_1235_58_n_1412));
  MX2X1 sub_1235_38_Y_add_1235_58_g2899(.A (instr_sub), .B
       (sub_1235_38_Y_add_1235_58_n_1443), .S0 (\reg_op2[2]_9671 ), .Y
       (sub_1235_38_Y_add_1235_58_n_1413));
  MX2X1 sub_1235_38_Y_add_1235_58_g2900(.A (instr_sub), .B
       (sub_1235_38_Y_add_1235_58_n_1443), .S0 (\reg_op2[19]_9688 ), .Y
       (sub_1235_38_Y_add_1235_58_n_1414));
  MX2X1 sub_1235_38_Y_add_1235_58_g2901(.A (instr_sub), .B
       (sub_1235_38_Y_add_1235_58_n_1443), .S0 (\reg_op2[7]_9676 ), .Y
       (sub_1235_38_Y_add_1235_58_n_1415));
  MX2X1 sub_1235_38_Y_add_1235_58_g2902(.A (instr_sub), .B
       (sub_1235_38_Y_add_1235_58_n_1443), .S0 (\reg_op2[24]_9693 ), .Y
       (sub_1235_38_Y_add_1235_58_n_1416));
  MX2X1 sub_1235_38_Y_add_1235_58_g2903(.A (instr_sub), .B
       (sub_1235_38_Y_add_1235_58_n_1443), .S0 (\reg_op2[1]_9670 ), .Y
       (sub_1235_38_Y_add_1235_58_n_1417));
  MX2X1 sub_1235_38_Y_add_1235_58_g2904(.A (instr_sub), .B
       (sub_1235_38_Y_add_1235_58_n_1443), .S0 (\reg_op2[16]_9685 ), .Y
       (sub_1235_38_Y_add_1235_58_n_1418));
  MX2X1 sub_1235_38_Y_add_1235_58_g2905(.A (instr_sub), .B
       (sub_1235_38_Y_add_1235_58_n_1443), .S0 (\reg_op2[9]_9678 ), .Y
       (sub_1235_38_Y_add_1235_58_n_1419));
  MX2X1 sub_1235_38_Y_add_1235_58_g2906(.A (instr_sub), .B
       (sub_1235_38_Y_add_1235_58_n_1443), .S0 (\reg_op2[20]_9689 ), .Y
       (sub_1235_38_Y_add_1235_58_n_1420));
  MX2X1 sub_1235_38_Y_add_1235_58_g2907(.A (instr_sub), .B
       (sub_1235_38_Y_add_1235_58_n_1443), .S0 (\reg_op2[21]_9690 ), .Y
       (sub_1235_38_Y_add_1235_58_n_1421));
  MX2X1 sub_1235_38_Y_add_1235_58_g2908(.A (instr_sub), .B
       (sub_1235_38_Y_add_1235_58_n_1443), .S0 (\reg_op2[3]_9672 ), .Y
       (sub_1235_38_Y_add_1235_58_n_1422));
  MX2X1 sub_1235_38_Y_add_1235_58_g2909(.A (instr_sub), .B
       (sub_1235_38_Y_add_1235_58_n_1443), .S0 (\reg_op2[26]_9695 ), .Y
       (sub_1235_38_Y_add_1235_58_n_1423));
  MX2X1 sub_1235_38_Y_add_1235_58_g2910(.A (instr_sub), .B
       (sub_1235_38_Y_add_1235_58_n_1443), .S0 (\reg_op2[14]_9683 ), .Y
       (sub_1235_38_Y_add_1235_58_n_1424));
  MX2X1 sub_1235_38_Y_add_1235_58_g2911(.A (instr_sub), .B
       (sub_1235_38_Y_add_1235_58_n_1443), .S0 (\reg_op2[0]_9669 ), .Y
       (sub_1235_38_Y_add_1235_58_n_1425));
  XNOR2X1 sub_1235_38_Y_add_1235_58_g2912(.A (\reg_op2[4]_9673 ), .B
       (sub_1235_38_Y_add_1235_58_n_1443), .Y
       (sub_1235_38_Y_add_1235_58_n_1426));
  XNOR2X1 sub_1235_38_Y_add_1235_58_g2913(.A (\reg_op2[22]_9691 ), .B
       (sub_1235_38_Y_add_1235_58_n_1443), .Y
       (sub_1235_38_Y_add_1235_58_n_1427));
  XNOR2X1 sub_1235_38_Y_add_1235_58_g2914(.A (\reg_op2[12]_9681 ), .B
       (sub_1235_38_Y_add_1235_58_n_1443), .Y
       (sub_1235_38_Y_add_1235_58_n_1428));
  XNOR2X1 sub_1235_38_Y_add_1235_58_g2915(.A (\reg_op2[11]_9680 ), .B
       (sub_1235_38_Y_add_1235_58_n_1443), .Y
       (sub_1235_38_Y_add_1235_58_n_1429));
  XNOR2X1 sub_1235_38_Y_add_1235_58_g2916(.A (\reg_op2[31]_9700 ), .B
       (sub_1235_38_Y_add_1235_58_n_1443), .Y
       (sub_1235_38_Y_add_1235_58_n_1430));
  XNOR2X1 sub_1235_38_Y_add_1235_58_g2917(.A (\reg_op2[29]_9698 ), .B
       (sub_1235_38_Y_add_1235_58_n_1443), .Y
       (sub_1235_38_Y_add_1235_58_n_1431));
  XNOR2X1 sub_1235_38_Y_add_1235_58_g2918(.A (\reg_op2[15]_9684 ), .B
       (sub_1235_38_Y_add_1235_58_n_1443), .Y
       (sub_1235_38_Y_add_1235_58_n_1432));
  XNOR2X1 sub_1235_38_Y_add_1235_58_g2919(.A (\reg_op2[17]_9686 ), .B
       (sub_1235_38_Y_add_1235_58_n_1443), .Y
       (sub_1235_38_Y_add_1235_58_n_1433));
  XNOR2X1 sub_1235_38_Y_add_1235_58_g2920(.A (\reg_op2[23]_9692 ), .B
       (sub_1235_38_Y_add_1235_58_n_1443), .Y
       (sub_1235_38_Y_add_1235_58_n_1434));
  XNOR2X1 sub_1235_38_Y_add_1235_58_g2921(.A (\reg_op2[8]_9677 ), .B
       (sub_1235_38_Y_add_1235_58_n_1443), .Y
       (sub_1235_38_Y_add_1235_58_n_1435));
  XNOR2X1 sub_1235_38_Y_add_1235_58_g2922(.A (\reg_op2[6]_9675 ), .B
       (sub_1235_38_Y_add_1235_58_n_1443), .Y
       (sub_1235_38_Y_add_1235_58_n_1436));
  XNOR2X1 sub_1235_38_Y_add_1235_58_g2923(.A (\reg_op2[30]_9699 ), .B
       (sub_1235_38_Y_add_1235_58_n_1443), .Y
       (sub_1235_38_Y_add_1235_58_n_1437));
  XNOR2X1 sub_1235_38_Y_add_1235_58_g2924(.A (\reg_op2[5]_9674 ), .B
       (sub_1235_38_Y_add_1235_58_n_1443), .Y
       (sub_1235_38_Y_add_1235_58_n_1438));
  XNOR2X1 sub_1235_38_Y_add_1235_58_g2925(.A (\reg_op2[25]_9694 ), .B
       (sub_1235_38_Y_add_1235_58_n_1443), .Y
       (sub_1235_38_Y_add_1235_58_n_1439));
  XNOR2X1 sub_1235_38_Y_add_1235_58_g2926(.A (\reg_op2[18]_9687 ), .B
       (sub_1235_38_Y_add_1235_58_n_1443), .Y
       (sub_1235_38_Y_add_1235_58_n_1440));
  XNOR2X1 sub_1235_38_Y_add_1235_58_g2927(.A (\reg_op2[13]_9682 ), .B
       (sub_1235_38_Y_add_1235_58_n_1443), .Y
       (sub_1235_38_Y_add_1235_58_n_1441));
  CLKXOR2X1 \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_g2492 (.A
       (n_7147), .B
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1132 ), .Y
       (\genblk2.pcpi_div_n_1930 ));
  ADDFX1 \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_g2493 (.A
       (\genblk2.pcpi_div_n_1867 ), .B (n_11719), .CI
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1134 ), .CO
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1132 ), .S
       (\genblk2.pcpi_div_n_1931 ));
  ADDFX1 \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_g2494 (.A
       (\genblk2.pcpi_div_n_1868 ), .B (n_11720), .CI
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1136 ), .CO
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1134 ), .S
       (\genblk2.pcpi_div_n_1932 ));
  ADDFX1 \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_g2495 (.A
       (\genblk2.pcpi_div_n_1869 ), .B (n_11729), .CI
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1138 ), .CO
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1136 ), .S
       (\genblk2.pcpi_div_n_1933 ));
  ADDFX1 \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_g2496 (.A
       (\genblk2.pcpi_div_n_1870 ), .B (n_11733), .CI
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1140 ), .CO
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1138 ), .S
       (\genblk2.pcpi_div_n_1934 ));
  ADDFX1 \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_g2497 (.A
       (\genblk2.pcpi_div_n_1871 ), .B (n_11722), .CI
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1142 ), .CO
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1140 ), .S
       (\genblk2.pcpi_div_n_1935 ));
  ADDFX1 \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_g2498 (.A
       (\genblk2.pcpi_div_n_1872 ), .B (n_11727), .CI
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1144 ), .CO
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1142 ), .S
       (\genblk2.pcpi_div_n_1936 ));
  ADDFX1 \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_g2499 (.A
       (\genblk2.pcpi_div_n_1873 ), .B (n_11714), .CI
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1146 ), .CO
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1144 ), .S
       (\genblk2.pcpi_div_n_1937 ));
  ADDFX1 \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_g2500 (.A
       (\genblk2.pcpi_div_n_1874 ), .B (n_11725), .CI
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1148 ), .CO
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1146 ), .S
       (\genblk2.pcpi_div_n_1938 ));
  ADDFX1 \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_g2501 (.A
       (\genblk2.pcpi_div_n_1875 ), .B (n_11726), .CI
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1150 ), .CO
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1148 ), .S
       (\genblk2.pcpi_div_n_1939 ));
  ADDFX1 \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_g2502 (.A
       (\genblk2.pcpi_div_n_1876 ), .B (n_11721), .CI
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1152 ), .CO
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1150 ), .S
       (\genblk2.pcpi_div_n_1940 ));
  ADDFX1 \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_g2503 (.A
       (\genblk2.pcpi_div_n_1877 ), .B (n_11706), .CI
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1154 ), .CO
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1152 ), .S
       (\genblk2.pcpi_div_n_1941 ));
  ADDFX1 \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_g2504 (.A
       (\genblk2.pcpi_div_n_1878 ), .B (n_11731), .CI
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1156 ), .CO
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1154 ), .S
       (\genblk2.pcpi_div_n_1942 ));
  ADDFX1 \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_g2505 (.A
       (\genblk2.pcpi_div_n_1879 ), .B (n_11723), .CI
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1158 ), .CO
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1156 ), .S
       (\genblk2.pcpi_div_n_1943 ));
  ADDFX1 \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_g2506 (.A
       (\genblk2.pcpi_div_n_1880 ), .B (n_11735), .CI
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1160 ), .CO
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1158 ), .S
       (\genblk2.pcpi_div_n_1944 ));
  ADDFX1 \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_g2507 (.A
       (\genblk2.pcpi_div_n_1881 ), .B (n_11715), .CI
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1162 ), .CO
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1160 ), .S
       (\genblk2.pcpi_div_n_1945 ));
  ADDFX1 \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_g2508 (.A
       (\genblk2.pcpi_div_n_1882 ), .B (n_11712), .CI
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1164 ), .CO
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1162 ), .S
       (\genblk2.pcpi_div_n_1946 ));
  ADDFX1 \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_g2509 (.A
       (\genblk2.pcpi_div_n_1883 ), .B (n_11711), .CI
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1166 ), .CO
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1164 ), .S
       (\genblk2.pcpi_div_n_1947 ));
  ADDFX1 \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_g2510 (.A
       (\genblk2.pcpi_div_n_1884 ), .B (n_11707), .CI
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1168 ), .CO
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1166 ), .S
       (\genblk2.pcpi_div_n_1948 ));
  ADDFX1 \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_g2511 (.A
       (\genblk2.pcpi_div_n_1885 ), .B (n_11732), .CI
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1170 ), .CO
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1168 ), .S
       (\genblk2.pcpi_div_n_1949 ));
  ADDFX1 \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_g2512 (.A
       (\genblk2.pcpi_div_n_1886 ), .B (n_11728), .CI
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1172 ), .CO
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1170 ), .S
       (\genblk2.pcpi_div_n_1950 ));
  ADDFX1 \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_g2513 (.A
       (\genblk2.pcpi_div_n_1887 ), .B (n_11718), .CI
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1174 ), .CO
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1172 ), .S
       (\genblk2.pcpi_div_n_1951 ));
  ADDFX1 \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_g2514 (.A
       (\genblk2.pcpi_div_n_1888 ), .B (n_11708), .CI
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1176 ), .CO
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1174 ), .S
       (\genblk2.pcpi_div_n_1952 ));
  ADDFX1 \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_g2515 (.A
       (\genblk2.pcpi_div_n_1889 ), .B (n_11734), .CI
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1178 ), .CO
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1176 ), .S
       (\genblk2.pcpi_div_n_1953 ));
  ADDFX1 \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_g2516 (.A
       (\genblk2.pcpi_div_n_1890 ), .B (n_11710), .CI
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1180 ), .CO
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1178 ), .S
       (\genblk2.pcpi_div_n_1954 ));
  ADDFX1 \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_g2517 (.A
       (\genblk2.pcpi_div_n_1891 ), .B (n_11730), .CI
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1182 ), .CO
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1180 ), .S
       (\genblk2.pcpi_div_n_1955 ));
  ADDFX1 \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_g2518 (.A
       (\genblk2.pcpi_div_n_1892 ), .B (n_11716), .CI
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1184 ), .CO
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1182 ), .S
       (\genblk2.pcpi_div_n_1956 ));
  ADDFX1 \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_g2519 (.A
       (\genblk2.pcpi_div_n_1893 ), .B (n_11724), .CI
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1186 ), .CO
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1184 ), .S
       (\genblk2.pcpi_div_n_1957 ));
  ADDFX1 \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_g2520 (.A
       (\genblk2.pcpi_div_n_1894 ), .B (n_11717), .CI
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1188 ), .CO
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1186 ), .S
       (\genblk2.pcpi_div_n_1958 ));
  ADDFX1 \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_g2521 (.A
       (\genblk2.pcpi_div_n_1895 ), .B (n_11713), .CI
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1190 ), .CO
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1188 ), .S
       (\genblk2.pcpi_div_n_1959 ));
  ADDFX1 \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_g2522 (.A
       (\genblk2.pcpi_div_n_1896 ), .B (n_11709), .CI
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1194 ), .CO
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1190 ), .S
       (\genblk2.pcpi_div_n_1960 ));
  OAI2BB1X1 \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_g2523 (.A0N
       (\genblk2.pcpi_div_n_1897 ), .A1N
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1213 ), .B0
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1194 ), .Y
       (\genblk2.pcpi_div_n_1961 ));
  NAND2BX1 \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_g2525 (.AN
       (\genblk2.pcpi_div_n_1897 ), .B (\genblk2.pcpi_div_n_1929 ), .Y
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1194 ));
  INVX1 \genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_g2543 (.A
       (\genblk2.pcpi_div_n_1929 ), .Y
       (\genblk2.pcpi_div_sub_2494_26_Y_minus_2469_59_n_1213 ));
  ADDFX1 add_1312_30_cdnfadd_2(.A (reg_pc[2]), .B (add_1312_30_n_1020),
       .CI (add_1312_30_n_991), .CO (add_1312_30_n_102), .S (n_6679));
  XNOR2X1 add_1312_30_g1255(.A (reg_pc[31]), .B (add_1312_30_n_851), .Y
       (n_6708));
  OA21X1 add_1312_30_g1256(.A0 (reg_pc[30]), .A1 (add_1312_30_n_856),
       .B0 (add_1312_30_n_851), .Y (n_6707));
  NAND2X1 add_1312_30_g1257(.A (reg_pc[30]), .B (add_1312_30_n_856), .Y
       (add_1312_30_n_851));
  AOI2BB1X1 add_1312_30_g1258(.A0N (reg_pc[29]), .A1N
       (add_1312_30_n_861), .B0 (add_1312_30_n_856), .Y (n_6706));
  AND2X1 add_1312_30_g1259(.A (add_1312_30_n_861), .B (reg_pc[29]), .Y
       (add_1312_30_n_856));
  AOI2BB1X1 add_1312_30_g1260(.A0N (reg_pc[28]), .A1N
       (add_1312_30_n_866), .B0 (add_1312_30_n_861), .Y (n_6705));
  AND2X1 add_1312_30_g1261(.A (add_1312_30_n_866), .B (reg_pc[28]), .Y
       (add_1312_30_n_861));
  AOI2BB1X1 add_1312_30_g1262(.A0N (reg_pc[27]), .A1N
       (add_1312_30_n_871), .B0 (add_1312_30_n_866), .Y (n_6704));
  AND2X1 add_1312_30_g1263(.A (add_1312_30_n_871), .B (reg_pc[27]), .Y
       (add_1312_30_n_866));
  AOI2BB1X1 add_1312_30_g1264(.A0N (reg_pc[26]), .A1N
       (add_1312_30_n_876), .B0 (add_1312_30_n_871), .Y (n_6703));
  AND2X1 add_1312_30_g1265(.A (add_1312_30_n_876), .B (reg_pc[26]), .Y
       (add_1312_30_n_871));
  AOI2BB1X1 add_1312_30_g1266(.A0N (reg_pc[25]), .A1N
       (add_1312_30_n_881), .B0 (add_1312_30_n_876), .Y (n_6702));
  AND2X1 add_1312_30_g1267(.A (add_1312_30_n_881), .B (reg_pc[25]), .Y
       (add_1312_30_n_876));
  AOI2BB1X1 add_1312_30_g1268(.A0N (reg_pc[24]), .A1N
       (add_1312_30_n_886), .B0 (add_1312_30_n_881), .Y (n_6701));
  AND2X1 add_1312_30_g1269(.A (add_1312_30_n_886), .B (reg_pc[24]), .Y
       (add_1312_30_n_881));
  AOI2BB1X1 add_1312_30_g1270(.A0N (reg_pc[23]), .A1N
       (add_1312_30_n_891), .B0 (add_1312_30_n_886), .Y (n_6700));
  AND2X1 add_1312_30_g1271(.A (add_1312_30_n_891), .B (reg_pc[23]), .Y
       (add_1312_30_n_886));
  AOI2BB1X1 add_1312_30_g1272(.A0N (reg_pc[22]), .A1N
       (add_1312_30_n_896), .B0 (add_1312_30_n_891), .Y (n_6699));
  AND2X1 add_1312_30_g1273(.A (add_1312_30_n_896), .B (reg_pc[22]), .Y
       (add_1312_30_n_891));
  AOI2BB1X1 add_1312_30_g1274(.A0N (reg_pc[21]), .A1N
       (add_1312_30_n_901), .B0 (add_1312_30_n_896), .Y (n_6698));
  AND2X1 add_1312_30_g1275(.A (add_1312_30_n_901), .B (reg_pc[21]), .Y
       (add_1312_30_n_896));
  AOI2BB1X1 add_1312_30_g1276(.A0N (reg_pc[20]), .A1N
       (add_1312_30_n_906), .B0 (add_1312_30_n_901), .Y (n_6697));
  AND2X1 add_1312_30_g1277(.A (add_1312_30_n_906), .B (reg_pc[20]), .Y
       (add_1312_30_n_901));
  AOI2BB1X1 add_1312_30_g1278(.A0N (reg_pc[19]), .A1N
       (add_1312_30_n_911), .B0 (add_1312_30_n_906), .Y (n_6696));
  AND2X1 add_1312_30_g1279(.A (add_1312_30_n_911), .B (reg_pc[19]), .Y
       (add_1312_30_n_906));
  AOI2BB1X1 add_1312_30_g1280(.A0N (reg_pc[18]), .A1N
       (add_1312_30_n_916), .B0 (add_1312_30_n_911), .Y (n_6695));
  AND2X1 add_1312_30_g1281(.A (add_1312_30_n_916), .B (reg_pc[18]), .Y
       (add_1312_30_n_911));
  AOI2BB1X1 add_1312_30_g1282(.A0N (reg_pc[17]), .A1N
       (add_1312_30_n_921), .B0 (add_1312_30_n_916), .Y (n_6694));
  AND2X1 add_1312_30_g1283(.A (add_1312_30_n_921), .B (reg_pc[17]), .Y
       (add_1312_30_n_916));
  AOI2BB1X1 add_1312_30_g1284(.A0N (reg_pc[16]), .A1N
       (add_1312_30_n_926), .B0 (add_1312_30_n_921), .Y (n_6693));
  AND2X1 add_1312_30_g1285(.A (add_1312_30_n_926), .B (reg_pc[16]), .Y
       (add_1312_30_n_921));
  AOI2BB1X1 add_1312_30_g1286(.A0N (reg_pc[15]), .A1N
       (add_1312_30_n_931), .B0 (add_1312_30_n_926), .Y (n_6692));
  AND2X1 add_1312_30_g1287(.A (add_1312_30_n_931), .B (reg_pc[15]), .Y
       (add_1312_30_n_926));
  AOI2BB1X1 add_1312_30_g1288(.A0N (reg_pc[14]), .A1N
       (add_1312_30_n_936), .B0 (add_1312_30_n_931), .Y (n_6691));
  AND2X1 add_1312_30_g1289(.A (add_1312_30_n_936), .B (reg_pc[14]), .Y
       (add_1312_30_n_931));
  AOI2BB1X1 add_1312_30_g1290(.A0N (reg_pc[13]), .A1N
       (add_1312_30_n_941), .B0 (add_1312_30_n_936), .Y (n_6690));
  AND2X1 add_1312_30_g1291(.A (add_1312_30_n_941), .B (reg_pc[13]), .Y
       (add_1312_30_n_936));
  AOI2BB1X1 add_1312_30_g1292(.A0N (reg_pc[12]), .A1N
       (add_1312_30_n_946), .B0 (add_1312_30_n_941), .Y (n_6689));
  AND2X1 add_1312_30_g1293(.A (add_1312_30_n_946), .B (reg_pc[12]), .Y
       (add_1312_30_n_941));
  AOI2BB1X1 add_1312_30_g1294(.A0N (reg_pc[11]), .A1N
       (add_1312_30_n_951), .B0 (add_1312_30_n_946), .Y (n_6688));
  AND2X1 add_1312_30_g1295(.A (add_1312_30_n_951), .B (reg_pc[11]), .Y
       (add_1312_30_n_946));
  AOI2BB1X1 add_1312_30_g1296(.A0N (reg_pc[10]), .A1N
       (add_1312_30_n_956), .B0 (add_1312_30_n_951), .Y (n_6687));
  AND2X1 add_1312_30_g1297(.A (add_1312_30_n_956), .B (reg_pc[10]), .Y
       (add_1312_30_n_951));
  AOI2BB1X1 add_1312_30_g1298(.A0N (reg_pc[9]), .A1N
       (add_1312_30_n_961), .B0 (add_1312_30_n_956), .Y (n_6686));
  AND2X1 add_1312_30_g1299(.A (add_1312_30_n_961), .B (reg_pc[9]), .Y
       (add_1312_30_n_956));
  AOI2BB1X1 add_1312_30_g1300(.A0N (reg_pc[8]), .A1N
       (add_1312_30_n_966), .B0 (add_1312_30_n_961), .Y (n_6685));
  AND2X1 add_1312_30_g1301(.A (add_1312_30_n_966), .B (reg_pc[8]), .Y
       (add_1312_30_n_961));
  AOI2BB1X1 add_1312_30_g1302(.A0N (reg_pc[7]), .A1N
       (add_1312_30_n_971), .B0 (add_1312_30_n_966), .Y (n_6684));
  AND2X1 add_1312_30_g1303(.A (add_1312_30_n_971), .B (reg_pc[7]), .Y
       (add_1312_30_n_966));
  AOI2BB1X1 add_1312_30_g1304(.A0N (reg_pc[6]), .A1N
       (add_1312_30_n_976), .B0 (add_1312_30_n_971), .Y (n_6683));
  AND2X1 add_1312_30_g1305(.A (add_1312_30_n_976), .B (reg_pc[6]), .Y
       (add_1312_30_n_971));
  AOI2BB1X1 add_1312_30_g1306(.A0N (reg_pc[5]), .A1N
       (add_1312_30_n_981), .B0 (add_1312_30_n_976), .Y (n_6682));
  AND2X1 add_1312_30_g1307(.A (add_1312_30_n_981), .B (reg_pc[5]), .Y
       (add_1312_30_n_976));
  AOI2BB1X1 add_1312_30_g1308(.A0N (reg_pc[4]), .A1N
       (add_1312_30_n_986), .B0 (add_1312_30_n_981), .Y (n_6681));
  AND2X1 add_1312_30_g1309(.A (add_1312_30_n_986), .B (reg_pc[4]), .Y
       (add_1312_30_n_981));
  AOI2BB1X1 add_1312_30_g1310(.A0N (reg_pc[3]), .A1N
       (add_1312_30_n_102), .B0 (add_1312_30_n_986), .Y (n_6680));
  AND2X1 add_1312_30_g1311(.A (add_1312_30_n_102), .B (reg_pc[3]), .Y
       (add_1312_30_n_986));
  ADDHX1 add_1312_30_g1312(.A (latched_compr), .B (reg_pc[1]), .CO
       (add_1312_30_n_991), .S (n_6678));
  INVX1 add_1312_30_g1313(.A (latched_compr), .Y (add_1312_30_n_1020));
  XNOR2X1 inc_add_382_74_g383(.A (n_6862), .B (inc_add_382_74_n_207),
       .Y (n_6832));
  NAND2X1 inc_add_382_74_g385(.A (n_6861), .B (inc_add_382_74_n_212),
       .Y (inc_add_382_74_n_207));
  NOR2BX1 inc_add_382_74_g387(.AN (n_6860), .B (inc_add_382_74_n_217),
       .Y (inc_add_382_74_n_212));
  NAND2X1 inc_add_382_74_g389(.A (n_6859), .B (inc_add_382_74_n_222),
       .Y (inc_add_382_74_n_217));
  AOI2BB1X1 inc_add_382_74_g390(.A0N (n_6858), .A1N
       (inc_add_382_74_n_227), .B0 (inc_add_382_74_n_222), .Y (n_6828));
  AND2X1 inc_add_382_74_g391(.A (inc_add_382_74_n_227), .B (n_6858), .Y
       (inc_add_382_74_n_222));
  AOI2BB1X1 inc_add_382_74_g392(.A0N (n_6857), .A1N
       (inc_add_382_74_n_232), .B0 (inc_add_382_74_n_227), .Y (n_6827));
  AND2X1 inc_add_382_74_g393(.A (inc_add_382_74_n_232), .B (n_6857), .Y
       (inc_add_382_74_n_227));
  NOR2BX1 inc_add_382_74_g395(.AN (n_6856), .B (inc_add_382_74_n_237),
       .Y (inc_add_382_74_n_232));
  NAND2X1 inc_add_382_74_g397(.A (n_6855), .B (inc_add_382_74_n_242),
       .Y (inc_add_382_74_n_237));
  AOI2BB1X1 inc_add_382_74_g398(.A0N (n_6854), .A1N
       (inc_add_382_74_n_247), .B0 (inc_add_382_74_n_242), .Y (n_6824));
  AND2X1 inc_add_382_74_g399(.A (inc_add_382_74_n_247), .B (n_6854), .Y
       (inc_add_382_74_n_242));
  NOR2BX1 inc_add_382_74_g401(.AN (n_6853), .B (inc_add_382_74_n_252),
       .Y (inc_add_382_74_n_247));
  NAND2X1 inc_add_382_74_g403(.A (n_6852), .B (inc_add_382_74_n_257),
       .Y (inc_add_382_74_n_252));
  AOI2BB1X1 inc_add_382_74_g404(.A0N (n_6851), .A1N
       (inc_add_382_74_n_262), .B0 (inc_add_382_74_n_257), .Y (n_6821));
  AND2X1 inc_add_382_74_g405(.A (inc_add_382_74_n_262), .B (n_6851), .Y
       (inc_add_382_74_n_257));
  NOR2BX1 inc_add_382_74_g407(.AN (n_6850), .B (inc_add_382_74_n_267),
       .Y (inc_add_382_74_n_262));
  XNOR2X1 inc_add_382_74_g408(.A (n_6849), .B (inc_add_382_74_n_272),
       .Y (n_6819));
  NAND2BX1 inc_add_382_74_g409(.AN (inc_add_382_74_n_272), .B (n_6849),
       .Y (inc_add_382_74_n_267));
  NAND2X1 inc_add_382_74_g411(.A (n_6848), .B (inc_add_382_74_n_277),
       .Y (inc_add_382_74_n_272));
  AOI2BB1X1 inc_add_382_74_g412(.A0N (n_6847), .A1N
       (inc_add_382_74_n_282), .B0 (inc_add_382_74_n_277), .Y (n_6817));
  AND2X1 inc_add_382_74_g413(.A (inc_add_382_74_n_282), .B (n_6847), .Y
       (inc_add_382_74_n_277));
  XNOR2X1 inc_add_382_74_g414(.A (n_6846), .B (inc_add_382_74_n_287),
       .Y (n_6816));
  NOR2BX1 inc_add_382_74_g415(.AN (n_6846), .B (inc_add_382_74_n_287),
       .Y (inc_add_382_74_n_282));
  OA21X1 inc_add_382_74_g416(.A0 (n_6845), .A1 (inc_add_382_74_n_292),
       .B0 (inc_add_382_74_n_287), .Y (n_6815));
  NAND2X1 inc_add_382_74_g417(.A (n_6845), .B (inc_add_382_74_n_292),
       .Y (inc_add_382_74_n_287));
  XNOR2X1 inc_add_382_74_g418(.A (n_6844), .B (inc_add_382_74_n_297),
       .Y (n_6814));
  NOR2BX1 inc_add_382_74_g419(.AN (n_6844), .B (inc_add_382_74_n_297),
       .Y (inc_add_382_74_n_292));
  OA21X1 inc_add_382_74_g420(.A0 (n_6843), .A1 (inc_add_382_74_n_302),
       .B0 (inc_add_382_74_n_297), .Y (n_6813));
  NAND2X1 inc_add_382_74_g421(.A (n_6843), .B (inc_add_382_74_n_302),
       .Y (inc_add_382_74_n_297));
  AOI2BB1X1 inc_add_382_74_g422(.A0N (n_6842), .A1N
       (inc_add_382_74_n_305), .B0 (inc_add_382_74_n_302), .Y (n_6812));
  AND2X1 inc_add_382_74_g423(.A (inc_add_382_74_n_305), .B (n_6842), .Y
       (inc_add_382_74_n_302));
  ADDHX1 inc_add_382_74_g424(.A (n_6841), .B (inc_add_382_74_n_309),
       .CO (inc_add_382_74_n_305), .S (n_6811));
  AOI2BB1X1 inc_add_382_74_g425(.A0N (n_6840), .A1N
       (inc_add_382_74_n_314), .B0 (inc_add_382_74_n_309), .Y (n_6810));
  AND2X1 inc_add_382_74_g426(.A (inc_add_382_74_n_314), .B (n_6840), .Y
       (inc_add_382_74_n_309));
  AOI2BB1X1 inc_add_382_74_g427(.A0N (n_6839), .A1N
       (inc_add_382_74_n_319), .B0 (inc_add_382_74_n_314), .Y (n_6809));
  AND2X1 inc_add_382_74_g428(.A (inc_add_382_74_n_319), .B (n_6839), .Y
       (inc_add_382_74_n_314));
  XNOR2X1 inc_add_382_74_g429(.A (n_6838), .B (inc_add_382_74_n_324),
       .Y (n_6808));
  NOR2BX1 inc_add_382_74_g430(.AN (n_6838), .B (inc_add_382_74_n_324),
       .Y (inc_add_382_74_n_319));
  OA21X1 inc_add_382_74_g431(.A0 (n_6837), .A1 (inc_add_382_74_n_329),
       .B0 (inc_add_382_74_n_324), .Y (n_6807));
  NAND2X1 inc_add_382_74_g432(.A (n_6837), .B (inc_add_382_74_n_329),
       .Y (inc_add_382_74_n_324));
  AOI2BB1X1 inc_add_382_74_g433(.A0N (n_6836), .A1N
       (inc_add_382_74_n_332), .B0 (inc_add_382_74_n_329), .Y (n_6806));
  AND2X1 inc_add_382_74_g434(.A (inc_add_382_74_n_332), .B (n_6836), .Y
       (inc_add_382_74_n_329));
  ADDHX1 inc_add_382_74_g435(.A (n_6835), .B (inc_add_382_74_n_336),
       .CO (inc_add_382_74_n_332), .S (n_6805));
  AOI2BB1X1 inc_add_382_74_g436(.A0N (n_6834), .A1N
       (inc_add_382_74_n_341), .B0 (inc_add_382_74_n_336), .Y (n_6804));
  AND2X1 inc_add_382_74_g437(.A (inc_add_382_74_n_341), .B (n_6834), .Y
       (inc_add_382_74_n_336));
  AOI2BB1X1 inc_add_382_74_g438(.A0N (n_6833), .A1N
       (mem_la_firstword_xfer), .B0 (inc_add_382_74_n_341), .Y
       (n_6803));
  AND2X1 inc_add_382_74_g439(.A (mem_la_firstword_xfer), .B (n_6833),
       .Y (inc_add_382_74_n_341));
  XNOR2X1 add_1864_26_g750(.A (add_1864_26_n_657), .B
       (add_1864_26_n_596), .Y (n_68));
  ADDFX1 add_1864_26_g751(.A (decoded_imm[30]), .B (\reg_op1[30]_9667
       ), .CI (add_1864_26_n_598), .CO (add_1864_26_n_596), .S (n_52));
  ADDFX1 add_1864_26_g752(.A (decoded_imm[29]), .B (\reg_op1[29]_9666
       ), .CI (add_1864_26_n_600), .CO (add_1864_26_n_598), .S
       (n_6931));
  ADDFX1 add_1864_26_g753(.A (decoded_imm[28]), .B (\reg_op1[28]_9665
       ), .CI (add_1864_26_n_602), .CO (add_1864_26_n_600), .S
       (n_6932));
  ADDFX1 add_1864_26_g754(.A (decoded_imm[27]), .B (\reg_op1[27]_9664
       ), .CI (add_1864_26_n_604), .CO (add_1864_26_n_602), .S
       (n_6933));
  ADDFX1 add_1864_26_g755(.A (decoded_imm[26]), .B (\reg_op1[26]_9663
       ), .CI (add_1864_26_n_606), .CO (add_1864_26_n_604), .S
       (n_6934));
  ADDFX1 add_1864_26_g756(.A (decoded_imm[25]), .B (\reg_op1[25]_9662
       ), .CI (add_1864_26_n_608), .CO (add_1864_26_n_606), .S
       (n_6935));
  ADDFX1 add_1864_26_g757(.A (decoded_imm[24]), .B (\reg_op1[24]_9661
       ), .CI (add_1864_26_n_610), .CO (add_1864_26_n_608), .S
       (n_6936));
  ADDFX1 add_1864_26_g758(.A (decoded_imm[23]), .B (\reg_op1[23]_9660
       ), .CI (add_1864_26_n_612), .CO (add_1864_26_n_610), .S
       (n_6937));
  ADDFX1 add_1864_26_g759(.A (decoded_imm[22]), .B (\reg_op1[22]_9659
       ), .CI (add_1864_26_n_614), .CO (add_1864_26_n_612), .S
       (n_6938));
  ADDFX1 add_1864_26_g760(.A (decoded_imm[21]), .B (\reg_op1[21]_9658
       ), .CI (add_1864_26_n_616), .CO (add_1864_26_n_614), .S
       (n_6939));
  ADDFX1 add_1864_26_g761(.A (decoded_imm[20]), .B (\reg_op1[20]_9657
       ), .CI (add_1864_26_n_618), .CO (add_1864_26_n_616), .S
       (n_6940));
  ADDFX1 add_1864_26_g762(.A (decoded_imm[19]), .B (\reg_op1[19]_9656
       ), .CI (add_1864_26_n_620), .CO (add_1864_26_n_618), .S
       (n_6941));
  ADDFX1 add_1864_26_g763(.A (decoded_imm[18]), .B (\reg_op1[18]_9655
       ), .CI (add_1864_26_n_622), .CO (add_1864_26_n_620), .S (n_50));
  ADDFX1 add_1864_26_g764(.A (decoded_imm[17]), .B (\reg_op1[17]_9654
       ), .CI (add_1864_26_n_624), .CO (add_1864_26_n_622), .S
       (n_6943));
  ADDFX1 add_1864_26_g765(.A (decoded_imm[16]), .B (\reg_op1[16]_9653
       ), .CI (add_1864_26_n_626), .CO (add_1864_26_n_624), .S
       (n_6944));
  ADDFX1 add_1864_26_g766(.A (decoded_imm[15]), .B (\reg_op1[15]_9652
       ), .CI (add_1864_26_n_628), .CO (add_1864_26_n_626), .S
       (n_6945));
  ADDFX1 add_1864_26_g767(.A (decoded_imm[14]), .B (\reg_op1[14]_9651
       ), .CI (add_1864_26_n_630), .CO (add_1864_26_n_628), .S (n_66));
  ADDFX1 add_1864_26_g768(.A (decoded_imm[13]), .B (\reg_op1[13]_9650
       ), .CI (add_1864_26_n_632), .CO (add_1864_26_n_630), .S
       (n_6947));
  ADDFX1 add_1864_26_g769(.A (decoded_imm[12]), .B (\reg_op1[12]_9649
       ), .CI (add_1864_26_n_634), .CO (add_1864_26_n_632), .S
       (n_6948));
  ADDFX1 add_1864_26_g770(.A (decoded_imm[11]), .B (\reg_op1[11]_9648
       ), .CI (add_1864_26_n_636), .CO (add_1864_26_n_634), .S
       (n_6949));
  ADDFX1 add_1864_26_g771(.A (decoded_imm[10]), .B (\reg_op1[10]_9647
       ), .CI (add_1864_26_n_638), .CO (add_1864_26_n_636), .S
       (n_6950));
  ADDFX1 add_1864_26_g772(.A (decoded_imm[9]), .B (\reg_op1[9]_9646 ),
       .CI (add_1864_26_n_640), .CO (add_1864_26_n_638), .S (n_6951));
  ADDFX1 add_1864_26_g773(.A (decoded_imm[8]), .B (\reg_op1[8]_9645 ),
       .CI (add_1864_26_n_642), .CO (add_1864_26_n_640), .S (n_6952));
  ADDFX1 add_1864_26_g774(.A (decoded_imm[7]), .B (\reg_op1[7]_9644 ),
       .CI (add_1864_26_n_644), .CO (add_1864_26_n_642), .S (n_6953));
  ADDFX1 add_1864_26_g775(.A (decoded_imm[6]), .B (\reg_op1[6]_9643 ),
       .CI (add_1864_26_n_646), .CO (add_1864_26_n_644), .S (n_6954));
  ADDFX1 add_1864_26_g776(.A (decoded_imm[5]), .B (\reg_op1[5]_9642 ),
       .CI (add_1864_26_n_648), .CO (add_1864_26_n_646), .S (n_6955));
  ADDFX1 add_1864_26_g777(.A (decoded_imm[4]), .B (\reg_op1[4]_9641 ),
       .CI (add_1864_26_n_650), .CO (add_1864_26_n_648), .S (n_6956));
  ADDFX1 add_1864_26_g778(.A (decoded_imm[3]), .B (\reg_op1[3]_9640 ),
       .CI (add_1864_26_n_652), .CO (add_1864_26_n_650), .S (n_114));
  ADDFX1 add_1864_26_g779(.A (decoded_imm[2]), .B (\reg_op1[2]_9639 ),
       .CI (add_1864_26_n_654), .CO (add_1864_26_n_652), .S (n_64));
  ADDFX1 add_1864_26_g780(.A (decoded_imm[1]), .B (\reg_op1[1]_9638 ),
       .CI (add_1864_26_n_658), .CO (add_1864_26_n_654), .S (n_62));
  AOI2BB1X1 add_1864_26_g781(.A0N (decoded_imm[0]), .A1N (reg_op1[0]),
       .B0 (add_1864_26_n_658), .Y (n_6960));
  XNOR2X1 add_1864_26_g782(.A (decoded_imm[31]), .B (\reg_op1[31]_9668
       ), .Y (add_1864_26_n_657));
  AND2X1 add_1864_26_g783(.A (reg_op1[0]), .B (decoded_imm[0]), .Y
       (add_1864_26_n_658));
  XNOR2X1 add_1801_23_g2358(.A (add_1801_23_n_1164), .B
       (add_1801_23_n_1105), .Y (n_115));
  ADDFX1 add_1801_23_g2359(.A (reg_pc[30]), .B (decoded_imm[30]), .CI
       (add_1801_23_n_1107), .CO (add_1801_23_n_1105), .S (n_112));
  ADDFX1 add_1801_23_g2360(.A (reg_pc[29]), .B (decoded_imm[29]), .CI
       (add_1801_23_n_1109), .CO (add_1801_23_n_1107), .S (n_110));
  ADDFX1 add_1801_23_g2361(.A (reg_pc[28]), .B (decoded_imm[28]), .CI
       (add_1801_23_n_1111), .CO (add_1801_23_n_1109), .S (n_106));
  ADDFX1 add_1801_23_g2362(.A (reg_pc[27]), .B (decoded_imm[27]), .CI
       (add_1801_23_n_1113), .CO (add_1801_23_n_1111), .S (n_108));
  ADDFX1 add_1801_23_g2363(.A (reg_pc[26]), .B (decoded_imm[26]), .CI
       (add_1801_23_n_1115), .CO (add_1801_23_n_1113), .S (n_104));
  ADDFX1 add_1801_23_g2364(.A (reg_pc[25]), .B (decoded_imm[25]), .CI
       (add_1801_23_n_1117), .CO (add_1801_23_n_1115), .S (n_102));
  ADDFX1 add_1801_23_g2365(.A (reg_pc[24]), .B (decoded_imm[24]), .CI
       (add_1801_23_n_1119), .CO (add_1801_23_n_1117), .S (n_100));
  ADDFX1 add_1801_23_g2366(.A (reg_pc[23]), .B (decoded_imm[23]), .CI
       (add_1801_23_n_1121), .CO (add_1801_23_n_1119), .S (n_98));
  ADDFX1 add_1801_23_g2367(.A (reg_pc[22]), .B (decoded_imm[22]), .CI
       (add_1801_23_n_1123), .CO (add_1801_23_n_1121), .S (n_96));
  ADDFX1 add_1801_23_g2368(.A (reg_pc[21]), .B (decoded_imm[21]), .CI
       (add_1801_23_n_1125), .CO (add_1801_23_n_1123), .S (n_94));
  ADDFX1 add_1801_23_g2369(.A (reg_pc[20]), .B (decoded_imm[20]), .CI
       (add_1801_23_n_1127), .CO (add_1801_23_n_1125), .S (n_88));
  ADDFX1 add_1801_23_g2370(.A (reg_pc[19]), .B (decoded_imm[19]), .CI
       (add_1801_23_n_1129), .CO (add_1801_23_n_1127), .S (n_92));
  ADDFX1 add_1801_23_g2371(.A (reg_pc[18]), .B (decoded_imm[18]), .CI
       (add_1801_23_n_1131), .CO (add_1801_23_n_1129), .S (n_90));
  ADDFX1 add_1801_23_g2372(.A (reg_pc[17]), .B (decoded_imm[17]), .CI
       (add_1801_23_n_1133), .CO (add_1801_23_n_1131), .S (n_86));
  ADDFX1 add_1801_23_g2373(.A (reg_pc[16]), .B (decoded_imm[16]), .CI
       (add_1801_23_n_1135), .CO (add_1801_23_n_1133), .S (n_6976));
  ADDFX1 add_1801_23_g2374(.A (reg_pc[15]), .B (decoded_imm[15]), .CI
       (add_1801_23_n_1137), .CO (add_1801_23_n_1135), .S (n_82));
  ADDFX1 add_1801_23_g2375(.A (reg_pc[14]), .B (decoded_imm[14]), .CI
       (add_1801_23_n_1139), .CO (add_1801_23_n_1137), .S (n_84));
  ADDFX1 add_1801_23_g2376(.A (reg_pc[13]), .B (decoded_imm[13]), .CI
       (add_1801_23_n_1141), .CO (add_1801_23_n_1139), .S (n_80));
  ADDFX1 add_1801_23_g2377(.A (reg_pc[12]), .B (decoded_imm[12]), .CI
       (add_1801_23_n_1143), .CO (add_1801_23_n_1141), .S (n_76));
  ADDFX1 add_1801_23_g2378(.A (reg_pc[11]), .B (decoded_imm[11]), .CI
       (add_1801_23_n_1145), .CO (add_1801_23_n_1143), .S (n_78));
  ADDFX1 add_1801_23_g2379(.A (reg_pc[10]), .B (decoded_imm[10]), .CI
       (add_1801_23_n_1147), .CO (add_1801_23_n_1145), .S (n_74));
  ADDFX1 add_1801_23_g2380(.A (reg_pc[9]), .B (decoded_imm[9]), .CI
       (add_1801_23_n_1149), .CO (add_1801_23_n_1147), .S (n_72));
  ADDFX1 add_1801_23_g2381(.A (reg_pc[8]), .B (decoded_imm[8]), .CI
       (add_1801_23_n_1151), .CO (add_1801_23_n_1149), .S (n_70));
  ADDFX1 add_1801_23_g2382(.A (reg_pc[7]), .B (decoded_imm[7]), .CI
       (add_1801_23_n_1153), .CO (add_1801_23_n_1151), .S (n_6985));
  ADDFX1 add_1801_23_g2383(.A (reg_pc[6]), .B (decoded_imm[6]), .CI
       (add_1801_23_n_1155), .CO (add_1801_23_n_1153), .S (n_6986));
  ADDFX1 add_1801_23_g2384(.A (reg_pc[5]), .B (decoded_imm[5]), .CI
       (add_1801_23_n_1157), .CO (add_1801_23_n_1155), .S (n_6987));
  ADDFX1 add_1801_23_g2385(.A (reg_pc[4]), .B (decoded_imm[4]), .CI
       (add_1801_23_n_1159), .CO (add_1801_23_n_1157), .S (n_6988));
  ADDFX1 add_1801_23_g2386(.A (reg_pc[3]), .B (decoded_imm[3]), .CI
       (add_1801_23_n_1161), .CO (add_1801_23_n_1159), .S (n_6989));
  ADDFX1 add_1801_23_g2387(.A (reg_pc[2]), .B (decoded_imm[2]), .CI
       (add_1801_23_n_1165), .CO (add_1801_23_n_1161), .S (n_6990));
  AOI2BB1X1 add_1801_23_g2388(.A0N (decoded_imm[1]), .A1N (reg_pc[1]),
       .B0 (add_1801_23_n_1165), .Y (n_54));
  XNOR2X1 add_1801_23_g2389(.A (reg_pc[31]), .B (decoded_imm[31]), .Y
       (add_1801_23_n_1164));
  AND2X1 add_1801_23_g2390(.A (decoded_imm[1]), .B (reg_pc[1]), .Y
       (add_1801_23_n_1165));
  XNOR2X1 add_1564_33_Y_add_1555_32_g732(.A
       (add_1564_33_Y_add_1555_32_n_645), .B
       (add_1564_33_Y_add_1555_32_n_585), .Y (n_6604));
  ADDFX1 add_1564_33_Y_add_1555_32_g733(.A (n_6624), .B
       (current_pc[30]), .CI (add_1564_33_Y_add_1555_32_n_587), .CO
       (add_1564_33_Y_add_1555_32_n_585), .S (n_6603));
  ADDFX1 add_1564_33_Y_add_1555_32_g734(.A (n_6624), .B
       (current_pc[29]), .CI (add_1564_33_Y_add_1555_32_n_590), .CO
       (add_1564_33_Y_add_1555_32_n_587), .S (n_6602));
  ADDFX1 add_1564_33_Y_add_1555_32_g735(.A (n_6624), .B
       (current_pc[28]), .CI (add_1564_33_Y_add_1555_32_n_592), .CO
       (add_1564_33_Y_add_1555_32_n_590), .S (n_6601));
  ADDFX1 add_1564_33_Y_add_1555_32_g736(.A (n_6624), .B
       (current_pc[27]), .CI (add_1564_33_Y_add_1555_32_n_594), .CO
       (add_1564_33_Y_add_1555_32_n_592), .S (n_6600));
  ADDFX1 add_1564_33_Y_add_1555_32_g737(.A (n_6624), .B
       (current_pc[26]), .CI (add_1564_33_Y_add_1555_32_n_596), .CO
       (add_1564_33_Y_add_1555_32_n_594), .S (n_6599));
  ADDFX1 add_1564_33_Y_add_1555_32_g738(.A (n_6624), .B
       (current_pc[25]), .CI (add_1564_33_Y_add_1555_32_n_598), .CO
       (add_1564_33_Y_add_1555_32_n_596), .S (n_6598));
  ADDFX1 add_1564_33_Y_add_1555_32_g739(.A (n_6624), .B
       (current_pc[24]), .CI (add_1564_33_Y_add_1555_32_n_600), .CO
       (add_1564_33_Y_add_1555_32_n_598), .S (n_6597));
  ADDFX1 add_1564_33_Y_add_1555_32_g740(.A (n_6624), .B
       (current_pc[23]), .CI (add_1564_33_Y_add_1555_32_n_602), .CO
       (add_1564_33_Y_add_1555_32_n_600), .S (n_6596));
  ADDFX1 add_1564_33_Y_add_1555_32_g741(.A (n_6624), .B
       (current_pc[22]), .CI (add_1564_33_Y_add_1555_32_n_604), .CO
       (add_1564_33_Y_add_1555_32_n_602), .S (n_6595));
  ADDFX1 add_1564_33_Y_add_1555_32_g742(.A (n_6624), .B
       (current_pc[21]), .CI (add_1564_33_Y_add_1555_32_n_606), .CO
       (add_1564_33_Y_add_1555_32_n_604), .S (n_6594));
  ADDFX1 add_1564_33_Y_add_1555_32_g743(.A (n_6624), .B
       (current_pc[20]), .CI (add_1564_33_Y_add_1555_32_n_608), .CO
       (add_1564_33_Y_add_1555_32_n_606), .S (n_6593));
  ADDFX1 add_1564_33_Y_add_1555_32_g744(.A (n_6623), .B
       (current_pc[19]), .CI (add_1564_33_Y_add_1555_32_n_610), .CO
       (add_1564_33_Y_add_1555_32_n_608), .S (n_6592));
  ADDFX1 add_1564_33_Y_add_1555_32_g745(.A (n_6622), .B
       (current_pc[18]), .CI (add_1564_33_Y_add_1555_32_n_612), .CO
       (add_1564_33_Y_add_1555_32_n_610), .S (n_6591));
  ADDFX1 add_1564_33_Y_add_1555_32_g746(.A (n_6621), .B
       (current_pc[17]), .CI (add_1564_33_Y_add_1555_32_n_614), .CO
       (add_1564_33_Y_add_1555_32_n_612), .S (n_6590));
  ADDFX1 add_1564_33_Y_add_1555_32_g747(.A (n_6620), .B
       (current_pc[16]), .CI (add_1564_33_Y_add_1555_32_n_616), .CO
       (add_1564_33_Y_add_1555_32_n_614), .S (n_6589));
  ADDFX1 add_1564_33_Y_add_1555_32_g748(.A (n_6619), .B
       (current_pc[15]), .CI (add_1564_33_Y_add_1555_32_n_618), .CO
       (add_1564_33_Y_add_1555_32_n_616), .S (n_6588));
  ADDFX1 add_1564_33_Y_add_1555_32_g749(.A (n_6618), .B
       (current_pc[14]), .CI (add_1564_33_Y_add_1555_32_n_620), .CO
       (add_1564_33_Y_add_1555_32_n_618), .S (n_6587));
  ADDFX1 add_1564_33_Y_add_1555_32_g750(.A (n_6617), .B
       (current_pc[13]), .CI (add_1564_33_Y_add_1555_32_n_622), .CO
       (add_1564_33_Y_add_1555_32_n_620), .S (n_6586));
  ADDFX1 add_1564_33_Y_add_1555_32_g751(.A (n_6616), .B
       (current_pc[12]), .CI (add_1564_33_Y_add_1555_32_n_624), .CO
       (add_1564_33_Y_add_1555_32_n_622), .S (n_6585));
  ADDFX1 add_1564_33_Y_add_1555_32_g752(.A (n_6615), .B
       (current_pc[11]), .CI (add_1564_33_Y_add_1555_32_n_626), .CO
       (add_1564_33_Y_add_1555_32_n_624), .S (n_6584));
  ADDFX1 add_1564_33_Y_add_1555_32_g753(.A (n_6614), .B
       (current_pc[10]), .CI (add_1564_33_Y_add_1555_32_n_628), .CO
       (add_1564_33_Y_add_1555_32_n_626), .S (n_6583));
  ADDFX1 add_1564_33_Y_add_1555_32_g754(.A (n_6613), .B
       (current_pc[9]), .CI (add_1564_33_Y_add_1555_32_n_630), .CO
       (add_1564_33_Y_add_1555_32_n_628), .S (n_6582));
  ADDFX1 add_1564_33_Y_add_1555_32_g755(.A (n_6612), .B
       (current_pc[8]), .CI (add_1564_33_Y_add_1555_32_n_632), .CO
       (add_1564_33_Y_add_1555_32_n_630), .S (n_6581));
  ADDFX1 add_1564_33_Y_add_1555_32_g756(.A (n_6611), .B
       (current_pc[7]), .CI (add_1564_33_Y_add_1555_32_n_634), .CO
       (add_1564_33_Y_add_1555_32_n_632), .S (n_6580));
  ADDFX1 add_1564_33_Y_add_1555_32_g757(.A (n_6610), .B
       (current_pc[6]), .CI (add_1564_33_Y_add_1555_32_n_636), .CO
       (add_1564_33_Y_add_1555_32_n_634), .S (n_6579));
  ADDFX1 add_1564_33_Y_add_1555_32_g758(.A (n_6609), .B
       (current_pc[5]), .CI (add_1564_33_Y_add_1555_32_n_638), .CO
       (add_1564_33_Y_add_1555_32_n_636), .S (n_6578));
  ADDFX1 add_1564_33_Y_add_1555_32_g759(.A (n_6608), .B
       (current_pc[4]), .CI (add_1564_33_Y_add_1555_32_n_640), .CO
       (add_1564_33_Y_add_1555_32_n_638), .S (n_6577));
  ADDFX1 add_1564_33_Y_add_1555_32_g760(.A (n_6607), .B
       (current_pc[3]), .CI (add_1564_33_Y_add_1555_32_n_642), .CO
       (add_1564_33_Y_add_1555_32_n_640), .S (n_6576));
  ADDFX1 add_1564_33_Y_add_1555_32_g761(.A (n_6606), .B
       (current_pc[2]), .CI (add_1564_33_Y_add_1555_32_n_646), .CO
       (add_1564_33_Y_add_1555_32_n_642), .S (n_6575));
  AOI2BB1X1 add_1564_33_Y_add_1555_32_g762(.A0N (n_6605), .A1N
       (current_pc[1]), .B0 (add_1564_33_Y_add_1555_32_n_646), .Y
       (n_6574));
  XNOR2X1 add_1564_33_Y_add_1555_32_g763(.A (n_6624), .B
       (current_pc[31]), .Y (add_1564_33_Y_add_1555_32_n_645));
  AND2X1 add_1564_33_Y_add_1555_32_g764(.A (current_pc[1]), .B
       (n_6605), .Y (add_1564_33_Y_add_1555_32_n_646));
  XNOR2X1 \genblk1.pcpi_mul_mul_2366_47_g47637 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1867 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2542 ), .Y
       (\genblk1.pcpi_mul_n_154 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47638 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1836 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1982 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2540 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2542 ), .S
       (\genblk1.pcpi_mul_n_153 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47639 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2056 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1983 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2538 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2540 ), .S
       (\genblk1.pcpi_mul_n_152 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47640 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2057 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2106 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2536 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2538 ), .S
       (\genblk1.pcpi_mul_n_151 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47641 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2107 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2144 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2534 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2536 ), .S
       (\genblk1.pcpi_mul_n_150 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47642 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2145 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2172 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2532 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2534 ), .S
       (\genblk1.pcpi_mul_n_149 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47643 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2238 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2173 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2530 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2532 ), .S
       (\genblk1.pcpi_mul_n_148 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47644 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2239 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2280 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2528 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2530 ), .S
       (\genblk1.pcpi_mul_n_147 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47645 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2288 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2281 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2526 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2528 ), .S
       (\genblk1.pcpi_mul_n_146 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47646 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2356 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2289 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2524 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2526 ), .S
       (\genblk1.pcpi_mul_n_145 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47647 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2357 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2338 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2522 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2524 ), .S
       (\genblk1.pcpi_mul_n_144 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47648 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2334 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2339 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2520 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2522 ), .S
       (\genblk1.pcpi_mul_n_143 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47649 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2344 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2335 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2518 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2520 ), .S
       (\genblk1.pcpi_mul_n_142 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47650 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2378 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2345 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2516 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2518 ), .S
       (\genblk1.pcpi_mul_n_141 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47651 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2364 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2379 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2514 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2516 ), .S
       (\genblk1.pcpi_mul_n_140 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47652 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2398 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2365 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2512 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2514 ), .S
       (\genblk1.pcpi_mul_n_139 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47653 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2404 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2399 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2510 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2512 ), .S
       (\genblk1.pcpi_mul_n_138 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47654 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2392 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2405 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2508 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2510 ), .S
       (\genblk1.pcpi_mul_n_137 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47655 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2406 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2393 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2506 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2508 ), .S
       (\genblk1.pcpi_mul_n_136 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47656 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2412 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2407 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2504 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2506 ), .S
       (\genblk1.pcpi_mul_n_135 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47657 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2414 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2413 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2502 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2504 ), .S
       (\genblk1.pcpi_mul_n_134 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47658 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2420 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2415 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2500 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2502 ), .S
       (\genblk1.pcpi_mul_n_133 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47659 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2422 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2421 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2498 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2500 ), .S
       (\genblk1.pcpi_mul_n_132 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47660 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2440 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2423 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2496 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2498 ), .S
       (\genblk1.pcpi_mul_n_131 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47661 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2438 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2441 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2494 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2496 ), .S
       (\genblk1.pcpi_mul_n_130 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47662 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2430 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2439 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2492 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2494 ), .S
       (\genblk1.pcpi_mul_n_129 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47663 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2428 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2431 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2490 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2492 ), .S
       (\genblk1.pcpi_mul_n_128 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47664 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2424 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2429 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2488 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2490 ), .S
       (\genblk1.pcpi_mul_n_127 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47665 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2432 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2425 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2486 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2488 ), .S
       (\genblk1.pcpi_mul_n_126 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47666 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2434 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2433 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2484 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2486 ), .S
       (\genblk1.pcpi_mul_n_125 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47667 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2418 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2435 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2482 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2484 ), .S
       (\genblk1.pcpi_mul_n_124 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47668 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2426 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2419 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2480 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2482 ), .S
       (\genblk1.pcpi_mul_n_123 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47669 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2416 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2427 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2478 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2480 ), .S
       (\genblk1.pcpi_mul_n_122 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47670 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2410 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2417 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2476 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2478 ), .S
       (\genblk1.pcpi_mul_n_121 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47671 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2402 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2411 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2474 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2476 ), .S
       (\genblk1.pcpi_mul_n_120 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47672 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2396 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2403 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2472 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2474 ), .S
       (\genblk1.pcpi_mul_n_119 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47673 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2384 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2397 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2470 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2472 ), .S
       (\genblk1.pcpi_mul_n_118 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47674 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2394 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2385 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2468 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2470 ), .S
       (\genblk1.pcpi_mul_n_117 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47675 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2400 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2395 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2466 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2468 ), .S
       (\genblk1.pcpi_mul_n_116 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47676 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2370 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2401 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2464 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2466 ), .S
       (\genblk1.pcpi_mul_n_115 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47677 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2360 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2371 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2462 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2464 ), .S
       (\genblk1.pcpi_mul_n_114 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47678 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2368 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2361 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2460 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2462 ), .S
       (\genblk1.pcpi_mul_n_113 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47679 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2342 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2369 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2458 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2460 ), .S
       (\genblk1.pcpi_mul_n_112 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47680 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2343 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2314 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2456 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2458 ), .S
       (\genblk1.pcpi_mul_n_111 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47681 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2312 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2315 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2454 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2456 ), .S
       (\genblk1.pcpi_mul_n_110 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47682 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2292 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2313 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2452 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2454 ), .S
       (\genblk1.pcpi_mul_n_109 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47683 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2293 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2268 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2450 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2452 ), .S
       (\genblk1.pcpi_mul_n_108 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47684 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2254 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2269 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2448 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2450 ), .S
       (\genblk1.pcpi_mul_n_107 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47685 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2272 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2255 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2446 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2448 ), .S
       (\genblk1.pcpi_mul_n_106 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47686 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2192 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2273 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2444 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2446 ), .S
       (\genblk1.pcpi_mul_n_105 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47687 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2132 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2193 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2442 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2444 ), .S
       (\genblk1.pcpi_mul_n_104 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47688 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2190 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2133 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2436 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2442 ), .S
       (\genblk1.pcpi_mul_n_103 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47689 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2318 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2387 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2382 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2440 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2441 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47690 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2286 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2383 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2366 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2438 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2439 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47691 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2090 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2191 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2408 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2436 ), .S
       (\genblk1.pcpi_mul_n_102 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47692 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2329 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2388 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2391 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2434 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2435 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47693 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2283 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2390 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2377 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2432 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2433 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47694 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2287 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2367 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2362 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2430 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2431 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47695 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2291 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2358 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2363 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2428 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2429 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47696 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2307 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2350 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2375 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2426 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2427 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47697 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2285 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2376 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2359 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2424 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2425 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47698 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2305 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2373 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2386 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2422 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2423 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47699 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2309 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2372 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2355 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2420 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2421 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47700 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2306 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2374 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2389 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2418 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2419 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47701 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2327 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2352 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2351 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2416 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2417 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47702 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2279 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2354 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2349 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2414 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2415 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47703 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2249 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2348 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2341 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2412 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2413 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47704 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2276 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2346 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2353 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2410 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2411 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47705 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2038 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2091 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2380 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2408 ), .S
       (\genblk1.pcpi_mul_n_101 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47706 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2185 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2340 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2311 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2406 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2407 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47707 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2155 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2317 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2294 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2404 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2405 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47708 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2277 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2332 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2347 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2402 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2403 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47709 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2153 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2296 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2321 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2400 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2401 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47710 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2165 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2301 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2316 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2398 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2399 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47711 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2215 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2322 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2333 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2396 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2397 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47712 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2161 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2320 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2299 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2394 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2395 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47713 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2184 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2310 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2295 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2392 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2393 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47714 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2266 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2247 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2336 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2390 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2391 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47715 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2183 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2267 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2337 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2388 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2389 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47716 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2234 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2163 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2325 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2386 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2387 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47717 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2237 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2298 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2323 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2384 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2385 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47718 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2230 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2235 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2319 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2382 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2383 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47719 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1872 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2039 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2330 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2380 ), .S
       (\genblk1.pcpi_mul_n_100 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47720 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2221 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2260 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2263 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2378 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2379 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47721 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2246 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2251 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2328 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2376 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2377 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47722 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2223 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2177 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2326 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2374 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2375 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47723 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2219 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2162 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2324 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2372 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2373 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47724 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2204 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2258 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2297 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2370 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2371 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47725 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2202 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2274 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2257 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2368 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2369 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47726 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2264 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2231 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2290 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2366 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2367 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47727 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2179 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2261 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2300 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2364 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2365 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47728 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2252 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2265 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2284 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2362 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2363 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47729 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2205 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2259 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2256 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2360 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2361 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47730 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2250 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2253 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2282 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2358 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2359 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47731 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1903 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2241 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2226 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2356 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2357 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47732 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2218 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2225 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2304 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2354 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2355 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47733 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2245 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2171 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2303 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2352 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2353 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47734 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2169 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2217 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2302 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2350 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2351 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47735 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2224 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2213 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2308 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2348 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2349 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47736 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2117 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2243 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2214 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2346 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2347 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47737 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2220 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2233 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2262 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2344 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2345 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47738 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2110 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2198 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2275 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2342 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2343 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47739 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2212 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2129 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2278 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2340 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2341 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47740 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2040 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2186 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2227 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2338 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2339 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47741 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2123 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2222 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2176 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2336 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2337 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47742 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2041 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2187 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2232 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2334 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2335 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47743 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2228 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2211 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2236 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2332 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2333 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47744 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1920 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1873 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2270 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2330 ), .S
       (\genblk1.pcpi_mul_n_99 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47745 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2182 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2125 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2127 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2328 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2329 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47746 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2013 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2244 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2170 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2326 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2327 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47747 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1980 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2167 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2158 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2324 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2325 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47748 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2208 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2229 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2160 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2322 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2323 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47749 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2112 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2157 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2150 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2320 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2321 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47750 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1981 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2206 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2159 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2318 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2319 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47751 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2180 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2115 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2200 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2316 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2317 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47752 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2111 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2196 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2199 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2314 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2315 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47753 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2087 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2194 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2197 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2312 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2313 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47754 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2128 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2109 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2248 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2310 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2311 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47755 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2007 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2119 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2174 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2308 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2309 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47756 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2121 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2168 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2216 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2306 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2307 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47757 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2079 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2175 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2166 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2304 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2305 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47758 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2116 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1997 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2242 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2302 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2303 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47759 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2114 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2071 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2154 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2300 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2301 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47760 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2156 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2209 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2152 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2298 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2299 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47761 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2034 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2113 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2151 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2296 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2297 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47762 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2108 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2181 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2201 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2294 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2295 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47763 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1943 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2142 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2195 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2292 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2293 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47764 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2137 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2140 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2139 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2290 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2291 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47765 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1875 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2240 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2103 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2288 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2289 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47766 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2136 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2138 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2207 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2286 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2287 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47767 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2134 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2130 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2141 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2284 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2285 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47768 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2124 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2135 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2131 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2282 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2283 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47769 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1874 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2101 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2102 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2280 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2281 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47770 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1923 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2105 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2118 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2278 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2279 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47771 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2005 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2066 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2210 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2276 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2277 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47772 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1959 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2021 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2203 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2274 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2275 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47773 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1935 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2044 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2095 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2272 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2273 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47774 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1839 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1921 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2188 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2270 ), .S
       (\genblk1.pcpi_mul_n_98 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47775 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2092 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2047 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2143 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2268 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2269 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47776 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1907 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2120 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1915 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2266 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2267 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47777 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1954 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2146 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1961 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2264 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2265 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47778 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2022 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1881 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2178 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2262 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2263 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47779 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2070 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2023 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2164 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2260 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2261 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47780 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2027 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2035 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2148 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2258 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2259 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47781 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2020 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2055 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2149 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2256 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2257 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47782 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2094 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1937 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2093 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2254 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2255 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47783 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1955 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1939 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2147 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2252 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2253 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47784 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1885 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1883 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2126 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2250 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2251 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47785 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2104 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1909 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2031 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2248 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2249 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47786 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1917 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2122 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1871 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2246 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2247 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47787 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1804 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2074 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2004 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2244 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2245 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47788 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1901 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2075 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1990 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2242 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2243 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47789 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1824 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2072 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1984 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2240 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2241 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47790 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2018 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2077 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2100 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2238 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2239 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47791 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2063 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2069 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2065 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2236 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2237 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47792 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2060 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1897 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2096 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2234 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2235 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47793 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1949 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1880 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2099 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2232 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2233 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47794 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1960 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2061 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2097 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2230 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2231 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47795 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1894 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1976 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1974 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2228 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2229 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47796 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2073 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1912 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1985 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2226 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2227 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47797 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2037 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2010 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2078 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2224 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2225 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47798 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1863 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1905 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2083 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2222 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2223 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47799 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1655 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2032 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1893 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2220 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2221 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47800 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2011 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2002 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1998 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2218 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2219 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47801 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2000 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2081 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2015 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2216 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2217 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47802 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2068 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1991 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2067 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2214 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2215 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47803 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1837 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1931 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2006 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2212 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2213 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47804 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2062 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2064 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1899 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2210 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2211 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47805 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1859 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1977 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1966 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2208 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2209 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47806 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1971 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1962 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1973 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2206 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2207 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47807 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2059 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2054 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1868 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2204 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2205 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47808 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1674 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1952 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2024 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2202 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2203 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47809 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2051 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2052 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1965 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2200 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2201 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47810 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1944 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2086 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2025 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2198 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2199 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47811 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2048 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1942 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1945 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2196 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2197 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47812 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1888 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2049 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2046 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2194 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2195 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47813 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1933 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2042 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2045 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2192 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2193 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47814 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1672 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1929 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1876 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2190 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2191 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47815 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1661 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1840 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2088 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2188 ), .S
       (\genblk1.pcpi_mul_n_97 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47816 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1913 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1948 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2098 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2186 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2187 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47817 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2030 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1908 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2053 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2184 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2185 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47818 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1904 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1911 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2028 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2182 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2183 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47819 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1780 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1857 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1926 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2180 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2181 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47820 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1841 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2008 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2033 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2178 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2179 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47821 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2014 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2012 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2029 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2176 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2177 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47822 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1613 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2016 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2085 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2174 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2175 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47823 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1843 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1879 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2076 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2172 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2173 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47824 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_2001 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1995 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1900 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2170 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2171 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47825 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1864 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1994 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1996 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2168 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2169 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47826 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1833 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1988 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2017 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2166 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2167 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47827 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1986 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2009 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1992 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2164 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2165 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47828 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1896 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2003 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1999 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2162 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2163 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47829 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1895 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1968 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1975 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2160 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2161 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47830 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1970 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1989 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1972 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2158 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2159 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47831 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1791 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1860 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1956 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2156 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2157 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47832 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1987 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1964 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1993 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2154 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2155 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47833 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1969 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1950 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1967 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2152 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2153 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47834 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1957 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_2026 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1951 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2150 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2151 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47835 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1958 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1856 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1869 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2148 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2149 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47836 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1853 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1830 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1946 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2146 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2147 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47837 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1637 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1891 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1878 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2144 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2145 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47838 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1827 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1889 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1936 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2142 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2143 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47839 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1882 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1884 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1941 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2140 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2141 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47840 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1963 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1979 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1938 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2138 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2139 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47841 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1718 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1829 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1940 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2136 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2137 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47842 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1849 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1924 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1947 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2134 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2135 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47843 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1852 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1928 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2043 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2132 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2133 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47844 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1854 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1916 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1870 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2130 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2131 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47845 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1930 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1922 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1887 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2128 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2129 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47846 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1850 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1914 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1925 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2126 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2127 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47847 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1647 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1910 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1906 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2124 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2125 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47848 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1648 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1786 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2082 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2122 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2123 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47849 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1682 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1620 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2080 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2120 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2121 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47850 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1540 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1838 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2084 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2118 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2119 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47851 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1796 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1861 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1898 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2116 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2117 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47852 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1779 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1594 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2050 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2114 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2115 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47853 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1798 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1792 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2058 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2112 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2113 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47854 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1516 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1865 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1953 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2110 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2111 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47855 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1858 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1886 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1927 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2108 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2109 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47856 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1560 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1846 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1890 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2106 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2107 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47857 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1646 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1514 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2036 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2104 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2105 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47858 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1746 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1823 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1902 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2102 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2103 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47859 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1745 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1574 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2019 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2100 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2101 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47860 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1694 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1832 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1892 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2098 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2099 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47861 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1717 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1568 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1978 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2096 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2097 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47862 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1680 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1628 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1932 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2094 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2095 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47863 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1679 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1828 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1934 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2092 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2093 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47864 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1480 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1847 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1877 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2090 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2091 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47865 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1535 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1662 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1918 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2088 ), .S
       (\genblk1.pcpi_mul_n_96 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47866 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1624 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1695 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1866 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2086 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2087 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47867 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1419 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1719 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1821 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2084 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2085 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47868 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1581 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1557 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1819 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2082 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2083 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47869 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1813 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1811 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1815 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2080 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2081 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47870 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1596 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1660 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1532 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2078 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2079 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47871 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1573 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1498 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1844 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2076 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2077 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47872 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1448 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1789 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1683 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2074 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2075 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47873 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1421 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1569 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1725 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2072 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2073 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47874 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1650 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1644 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1842 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2070 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2071 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47875 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1578 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1774 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1768 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2068 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2069 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47876 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1767 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1790 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1862 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2066 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2067 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47877 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1765 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1572 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1778 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2064 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2065 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47878 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1551 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1729 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1761 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2062 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2063 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47879 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1512 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1738 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1564 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2060 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2061 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47880 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1450 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1723 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1759 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2058 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2059 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47881 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1559 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1782 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1845 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2056 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2057 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47882 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1673 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1760 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1652 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2054 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2055 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47883 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1538 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1754 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1548 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2052 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2053 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47884 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1753 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1537 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1547 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2050 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2051 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47885 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1469 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1617 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1691 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2048 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2049 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47886 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1470 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1618 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1692 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2046 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2047 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47887 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1708 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1706 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1851 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2044 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2045 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47888 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1714 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1716 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1671 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2042 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2043 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47889 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1570 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1770 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1831 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2040 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2041 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47890 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1787 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1602 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1848 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2038 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2039 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47891 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1595 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1799 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1659 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2036 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2037 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47892 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1476 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1542 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1855 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2034 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2035 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47893 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1633 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1649 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1643 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2032 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2033 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47894 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1645 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1712 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1732 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2030 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2031 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47895 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1640 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1616 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1520 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2028 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2029 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47896 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1651 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1562 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1734 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2026 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2027 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47897 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1805 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1636 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1690 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2024 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2025 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47898 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1528 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1740 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1656 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2022 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2023 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47899 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1482 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1622 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1600 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2020 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2021 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47900 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1185 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1735 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1590 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2018 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2019 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47901 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1607 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1605 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1609 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2016 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2017 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47902 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1803 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1820 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1632 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2014 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2015 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47903 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1464 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1558 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1582 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2012 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2013 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47904 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1741 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1625 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1800 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2010 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2011 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47905 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1653 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1593 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1634 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2008 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2009 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47906 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1668 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1678 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1676 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2006 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2007 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47907 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1586 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1794 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1808 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2004 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2005 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47908 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1545 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1742 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1720 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2002 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2003 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47909 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1807 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1795 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1818 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_2000 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_2001 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47910 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1614 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1626 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1822 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1998 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1999 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47911 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1812 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1814 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1816 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1996 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1997 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47912 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1585 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1793 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1587 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1994 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1995 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47913 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1783 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1654 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1612 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1992 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1993 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47914 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1510 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1554 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1684 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1990 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1991 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47915 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1567 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1709 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1737 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1988 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1989 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47916 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1423 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1771 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1763 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1986 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1987 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47917 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1769 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1468 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1502 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1984 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1985 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47918 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1428 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1781 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1472 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1982 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1983 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47919 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1610 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1606 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1834 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1980 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1981 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47920 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1521 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1727 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1743 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1978 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1979 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47921 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1757 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1751 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1766 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1976 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1977 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47922 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1552 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1762 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1730 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1974 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1975 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47923 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1755 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1657 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1710 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1972 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1973 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47924 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1426 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1747 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1529 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1970 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1971 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47925 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1749 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1797 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1752 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1968 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1969 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47926 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1508 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1544 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1758 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1966 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1967 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47927 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1784 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1772 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1764 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1964 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1965 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47928 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1641 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1523 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1748 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1962 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1963 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47929 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1756 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1658 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1530 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1960 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1961 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47930 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1635 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1515 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1689 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1958 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1959 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47931 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1475 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1733 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1541 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1956 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1957 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47932 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1524 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1522 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1642 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1954 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1955 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47933 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1441 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1591 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1623 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1952 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1953 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47934 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1561 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1750 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1776 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1950 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1951 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47935 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1721 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1489 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1484 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1948 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1949 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47936 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1579 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1575 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1699 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1946 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1947 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47937 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1592 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1697 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1806 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1944 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1945 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47938 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1696 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1702 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1698 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1942 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1943 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47939 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1499 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1473 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1687 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1940 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1941 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47940 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1495 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1744 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1728 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1938 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1939 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47941 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1627 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1486 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1686 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1936 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1937 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47942 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1492 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1705 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1707 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1934 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1935 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47943 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1438 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1713 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1715 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1932 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1933 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47944 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1539 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1677 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1675 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1930 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1931 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47945 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1479 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1669 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1534 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1928 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1929 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47946 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1517 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1711 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1731 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1926 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1927 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47947 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1785 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1665 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1663 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1924 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1925 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47948 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1667 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1506 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1478 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1922 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1923 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47949 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1443 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1583 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1598 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1920 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1921 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47950 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1413 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1536 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1825 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1918 ), .S
       (\genblk1.pcpi_mul_n_95 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47951 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1809 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1550 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1466 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1916 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1917 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47952 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1666 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1810 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1664 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1914 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1915 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47953 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1693 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1483 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1726 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1912 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1913 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47954 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1519 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1566 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1681 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1910 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1911 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47955 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1513 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1518 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1704 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1908 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1909 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47956 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1639 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1615 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1619 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1906 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1907 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47957 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1444 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1463 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1631 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1904 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1905 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47958 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1501 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1504 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1488 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1902 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1903 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47959 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1553 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1509 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1588 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1900 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1901 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47960 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1571 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1773 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1577 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1898 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1899 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47961 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1511 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1546 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1608 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1896 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1897 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47962 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1459 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1507 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1543 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1894 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1895 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47963 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1187 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1527 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1739 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1892 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1893 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47964 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1178 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1493 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1802 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1890 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1891 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47965 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1314 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1485 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1685 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1888 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1889 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47966 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1183 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1477 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1505 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1886 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1887 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47967 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1465 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1496 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1688 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1884 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1885 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47968 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1474 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1556 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1500 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1882 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1883 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47969 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1722 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1490 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1526 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1880 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1881 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47970 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1497 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1494 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1638 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1878 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1879 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47971 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1446 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1601 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1670 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1876 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1877 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47972 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1503 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1487 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1736 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1874 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1875 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47973 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1597 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1604 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1788 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1872 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1873 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47974 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1700 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1580 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1576 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1870 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1871 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47975 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1481 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1599 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1724 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1868 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1869 ));
  XNOR2X1 \genblk1.pcpi_mul_mul_2366_47_g47976 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1462 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1835 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1867 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47977 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1011 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1332 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1701 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1865 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1866 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47978 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1248 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1279 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1817 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1863 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1864 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47979 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_990 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1458 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1777 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1861 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1862 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47980 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1216 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1449 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1775 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1859 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1860 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47981 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1017 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1190 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1703 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1857 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1858 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47982 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1049 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1455 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1621 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1855 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1856 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47983 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1180 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1453 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1549 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1853 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1854 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47984 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1018 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1447 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1533 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1851 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1852 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47985 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1063 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1565 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1461 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1849 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1850 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47986 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_932 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1603 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1454 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1847 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1848 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47987 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1243 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1177 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1801 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1845 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1846 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47988 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_977 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1425 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1589 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1843 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1844 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47989 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1422 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1200 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1611 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1841 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1842 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47990 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1326 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1323 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1584 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1839 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1840 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47991 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1241 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1418 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1531 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1837 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1838 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47992 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_881 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1232 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1471 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1835 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1836 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47993 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_969 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1417 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1563 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1833 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1834 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47994 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1213 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1182 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1525 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1831 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1832 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47995 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1203 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1179 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1555 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1829 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1830 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47996 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1310 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1439 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1491 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1827 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1828 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47997 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1414 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1445 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1629 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1825 ), .S
       (\genblk1.pcpi_mul_n_94 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47998 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_909 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1420 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1467 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1823 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1824 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g47999 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1246 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1358 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1249 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1821 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1822 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48000 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1042 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1130 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1278 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1819 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1820 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48001 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1247 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1359 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1319 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1817 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1818 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48002 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1367 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1265 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1264 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1815 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1816 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48003 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1262 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1365 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1260 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1813 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1814 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48004 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1258 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1257 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1363 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1811 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1812 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48005 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1313 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1308 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1391 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1809 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1810 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48006 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1215 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1214 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1344 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1807 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1808 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48007 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1014 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1380 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1013 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1805 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1806 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48008 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1357 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1242 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1442 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1803 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1804 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48009 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_873 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1400 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1045 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1801 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1802 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48010 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_860 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1297 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1382 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1799 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1800 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48011 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1065 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1097 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1066 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1797 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1798 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48012 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1343 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1211 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1210 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1795 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1796 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48013 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_843 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1317 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1346 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1793 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1794 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48014 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1084 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1060 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1460 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1791 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1792 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48015 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1227 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1337 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1196 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1789 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1790 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48016 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1174 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1266 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1229 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1787 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1788 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48017 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1207 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1397 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_937 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1785 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1786 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48018 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_878 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1230 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1099 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1783 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1784 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48019 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_854 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1429 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_989 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1781 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1782 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48020 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1078 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1081 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1189 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1779 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1780 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48021 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_845 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1309 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1094 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1777 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1778 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48022 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1092 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1070 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1071 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1775 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1776 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48023 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_938 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1162 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_939 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1773 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1774 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48024 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1062 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_4 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1096 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1771 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1772 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48025 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1228 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1181 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1068 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1769 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1770 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48026 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1022 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_973 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1451 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1767 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1768 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48027 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_986 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1140 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_987 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1765 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1766 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48028 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1105 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1032 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1040 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1763 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1764 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48029 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_991 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1131 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1002 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1761 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1762 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48030 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1061 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1176 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1059 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1759 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1760 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48031 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_840 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1304 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1113 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1757 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1758 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48032 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1086 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1088 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1089 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1755 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1756 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48033 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1055 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1051 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1104 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1753 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1754 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48034 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1036 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1108 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1037 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1751 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1752 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48035 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_863 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1152 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1058 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1749 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1750 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48036 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1098 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1041 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1072 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1747 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1748 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48037 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_869 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_996 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1186 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1745 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1746 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48038 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_892 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1039 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1111 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1743 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1744 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48039 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1193 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_7 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1336 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1741 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1742 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48040 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_944 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1012 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1383 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1739 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1740 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48041 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1006 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1125 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_3 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1737 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1738 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48042 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1212 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1171 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1057 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1735 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1736 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48043 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1083 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1164 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1082 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1733 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1734 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48044 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1307 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1137 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1004 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1731 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1732 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48045 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1133 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1000 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1001 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1729 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1730 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48046 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1048 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1106 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_0 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1727 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1728 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48047 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1009 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1119 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_5 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1725 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1726 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48048 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_861 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1101 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1064 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1723 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1724 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48049 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_901 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1195 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1167 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1721 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1722 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48050 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1254 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1253 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1360 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1719 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1720 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48051 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_914 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1223 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1427 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1717 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1718 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48052 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_842 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1169 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1280 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1715 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1716 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48053 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_877 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1155 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_963 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1713 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1714 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48054 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1024 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_9 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1143 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1711 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1712 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48055 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1141 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_983 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_978 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1709 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1710 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48056 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1138 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_955 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_966 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1707 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1708 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48057 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1231 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1149 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1283 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1705 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1706 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48058 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1208 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1128 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1316 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1703 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1704 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48059 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_958 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1145 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1010 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1701 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1702 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48060 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_981 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_979 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1147 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1699 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1700 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48061 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1007 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1292 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1129 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1697 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1698 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48062 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1003 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1386 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1440 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1695 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1696 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48063 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_894 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_998 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1390 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1693 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1694 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48064 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_943 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1139 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_997 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1691 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1692 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48065 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1318 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1372 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1031 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1689 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1690 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48066 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_968 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_967 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1157 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1687 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1688 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48067 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_984 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1160 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_982 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1685 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1686 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48068 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1074 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1375 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1197 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1683 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1684 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48069 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1268 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1153 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1052 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1681 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1682 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48070 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1046 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1393 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1331 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1679 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1680 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48071 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1334 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1387 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1677 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1678 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48072 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1151 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1069 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1325 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1675 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1676 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48073 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1038 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1376 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1328 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1673 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1674 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48074 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1076 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_949 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1456 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1671 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1672 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48075 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_850 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1352 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1270 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1669 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1670 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48076 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1008 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1315 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1370 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1667 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1668 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48077 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_992 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1016 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1389 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1665 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1666 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48078 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1126 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_975 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1329 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1663 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1664 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48079 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1348 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1273 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1437 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1661 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1662 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48080 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1289 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1288 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1378 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1659 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1660 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48081 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1075 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1322 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1091 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1657 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1658 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48082 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1188 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1277 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1275 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1655 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1656 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48083 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_905 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1300 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1175 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1653 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1654 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48084 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1054 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1132 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1053 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1651 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1652 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48085 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1256 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_10 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1362 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1649 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1650 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48086 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_999 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1311 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1379 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1647 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1648 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48087 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_961 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1301 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1184 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1645 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1646 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48088 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1251 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1356 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1244 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1643 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1644 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48089 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1118 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_941 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1028 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1641 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1642 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48090 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1403 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1296 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1324 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1639 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1640 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48091 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_910 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1282 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1424 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1637 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1638 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48092 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_942 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1117 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1029 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1635 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1636 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48093 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_899 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1233 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1351 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1633 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1634 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48094 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1286 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1285 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1377 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1631 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1632 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48095 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_851 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_880 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1430 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1629 ), .S
       (\genblk1.pcpi_mul_n_93 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48096 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1035 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1148 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1015 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1627 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1628 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48097 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1238 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1234 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1364 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1625 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1626 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48098 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1050 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1124 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1293 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1623 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1624 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48099 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1047 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1107 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1299 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1621 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1622 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48100 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1303 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1361 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_948 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1619 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1620 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48101 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1142 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_994 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_993 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1617 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1618 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48102 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1295 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1294 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1381 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1615 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1616 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48103 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_908 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1416 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1349 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1613 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1614 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48104 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1245 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1338 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1194 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1611 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1612 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48105 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1392 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1222 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1224 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1609 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1610 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48106 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1219 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1217 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1345 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1607 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1608 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48107 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1206 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1209 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1340 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1605 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1606 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48108 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_848 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_867 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1384 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1603 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1604 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48109 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_874 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1136 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_934 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1601 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1602 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48110 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1116 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1298 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1033 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1599 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1600 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48111 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1396 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1333 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1335 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1597 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1598 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48112 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1255 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1291 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1412 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1595 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1596 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48113 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_936 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1161 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_933 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1593 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1594 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48114 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_846 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_855 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1121 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1591 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1592 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48115 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_898 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1402 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1026 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1589 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1590 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48116 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1239 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1347 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1226 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1587 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1588 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48117 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_868 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1220 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1395 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1585 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1586 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48118 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_839 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_858 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1411 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1583 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1584 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48119 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1271 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1272 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1371 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1581 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1582 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48120 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_821 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1287 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1388 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1579 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1580 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48121 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_945 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1158 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_947 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1577 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1578 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48122 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_950 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_959 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1144 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1575 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1576 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48123 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_13 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1166 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1034 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1573 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1574 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48124 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_857 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_935 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1168 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1571 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1572 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48125 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_912 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1281 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1374 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1569 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1570 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48126 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1134 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_951 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_995 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1567 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1568 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48127 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_911 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_871 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1404 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1565 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1566 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48128 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_970 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1394 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_964 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1563 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1564 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48129 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1330 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1095 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1073 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1561 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1562 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48130 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_895 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_12 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1366 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1559 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1560 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48131 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1276 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1274 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1373 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1557 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1558 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48132 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_906 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_988 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1406 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1555 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1556 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48133 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_866 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1205 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1341 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1553 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1554 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48134 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_865 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1005 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1127 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1551 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1552 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48135 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_915 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1204 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1135 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1549 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1550 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48136 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1103 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1056 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_960 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1547 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1548 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48137 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_900 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1235 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1165 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1545 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1546 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48138 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1021 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1115 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1025 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1543 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1544 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48139 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_838 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1087 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1407 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1541 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1542 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48140 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_913 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1263 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1114 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1539 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1540 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48141 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_893 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1221 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1110 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1537 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1538 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48142 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_844 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_876 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1410 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1535 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1536 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48143 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_853 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_954 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1159 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1533 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1534 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48144 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1354 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1240 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1077 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1531 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1532 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48145 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1080 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1079 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1093 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1529 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1530 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48146 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_862 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_940 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1399 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1527 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1528 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48147 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1027 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1350 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_2 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1525 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1526 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48148 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1023 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1019 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1123 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1523 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1524 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48149 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1044 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1043 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1122 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1521 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1522 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48150 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1306 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1305 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1369 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1519 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1520 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48151 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_902 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_985 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1154 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1517 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1518 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48152 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1172 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1030 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1320 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1515 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1516 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48153 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1259 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1385 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1067 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1513 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1514 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48154 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_896 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1261 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1102 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1511 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1512 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48155 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1202 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1339 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1201 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1509 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1510 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48156 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_864 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1120 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1020 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1507 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1508 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48157 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1170 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_953 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_956 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1505 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1506 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48158 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1267 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_11 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1302 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1503 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1504 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48159 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_904 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1237 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1173 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1501 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1502 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48160 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_972 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_971 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1150 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1499 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1500 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48161 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_907 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1401 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1198 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1497 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1498 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48162 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1199 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_962 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1100 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1495 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1496 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48163 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1250 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_8 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_976 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1493 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1494 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48164 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_849 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_870 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1408 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1491 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1492 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48165 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1109 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1327 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1321 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1489 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1490 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48166 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1252 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1368 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1269 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1487 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1488 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48167 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1146 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_980 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1284 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1485 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1486 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48168 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1398 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1290 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1236 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1483 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1484 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48169 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_837 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_859 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1112 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1481 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1482 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48170 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_875 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1163 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_946 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1479 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1480 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48171 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_903 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1312 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1355 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1477 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1478 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48172 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_852 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1085 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1090 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1475 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1476 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48173 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1353 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_974 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_952 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1473 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1474 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48174 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_897 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1192 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_6 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1471 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1472 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48175 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_841 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_856 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1405 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1469 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1470 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48176 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1218 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1342 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1225 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1467 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1468 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48177 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_957 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_965 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1156 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1465 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1466 ));
  ADDFX1 \genblk1.pcpi_mul_mul_2366_47_g48178 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_847 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_872 ), .CI
       (\genblk1.pcpi_mul_mul_2366_47_n_1409 ), .CO
       (\genblk1.pcpi_mul_mul_2366_47_n_1463 ), .S
       (\genblk1.pcpi_mul_mul_2366_47_n_1464 ));
  XNOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48179 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_881 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1457 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1462 ));
  OAI2BB1X1 \genblk1.pcpi_mul_mul_2366_47_g48180 (.A0N
       (\genblk1.pcpi_mul_mul_2366_47_n_931 ), .A1N
       (\genblk1.pcpi_mul_mul_2366_47_n_1191 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_1453 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1461 ));
  XNOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48181 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_919 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1432 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1460 ));
  XNOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48182 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_921 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1435 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1459 ));
  XNOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48183 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_920 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1436 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1458 ));
  XNOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48184 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_879 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1415 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1457 ));
  XNOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48185 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_916 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1433 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1456 ));
  XNOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48186 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_917 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1434 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1455 ));
  XNOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48187 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_923 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1431 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1454 ));
  AOI21X1 \genblk1.pcpi_mul_mul_2366_47_g48188 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_819 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_891 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_1430 ), .Y
       (\genblk1.pcpi_mul_n_92 ));
  NOR2BX1 \genblk1.pcpi_mul_mul_2366_47_g48189 (.AN
       (\genblk1.pcpi_mul_mul_2366_47_n_1435 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_921 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1451 ));
  NOR2BX1 \genblk1.pcpi_mul_mul_2366_47_g48190 (.AN
       (\genblk1.pcpi_mul_mul_2366_47_n_1434 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_917 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1450 ));
  NOR2BX1 \genblk1.pcpi_mul_mul_2366_47_g48191 (.AN
       (\genblk1.pcpi_mul_mul_2366_47_n_1432 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_919 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1449 ));
  NOR2BX1 \genblk1.pcpi_mul_mul_2366_47_g48192 (.AN
       (\genblk1.pcpi_mul_mul_2366_47_n_1436 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_920 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1448 ));
  NOR2BX1 \genblk1.pcpi_mul_mul_2366_47_g48193 (.AN
       (\genblk1.pcpi_mul_mul_2366_47_n_1433 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_916 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1447 ));
  NOR2BX1 \genblk1.pcpi_mul_mul_2366_47_g48194 (.AN
       (\genblk1.pcpi_mul_mul_2366_47_n_1431 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_923 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1446 ));
  OR2X1 \genblk1.pcpi_mul_mul_2366_47_g48195 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_931 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_1191 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1453 ));
  XNOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48196 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_927 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_890 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1445 ));
  XNOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48197 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_930 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_884 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1444 ));
  XNOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48198 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_922 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_883 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1443 ));
  XNOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48199 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_926 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_888 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1442 ));
  XNOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48200 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_918 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_885 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1441 ));
  XNOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48201 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_928 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_886 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1440 ));
  XNOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48202 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_925 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_882 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1439 ));
  XNOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48203 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_929 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_889 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1438 ));
  XNOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48204 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_924 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_887 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1437 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_g48205 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1428 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1429 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_g48206 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1426 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1427 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_g48207 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1424 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1425 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_g48208 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1422 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1423 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_g48209 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1420 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1421 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_g48210 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1418 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1419 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_g48211 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1416 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1417 ));
  AOI21X1 \genblk1.pcpi_mul_mul_2366_47_g48212 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_836 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_789 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1415 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48213 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_247 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_835 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_788 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1414 ));
  NOR2BX1 \genblk1.pcpi_mul_mul_2366_47_g48214 (.AN
       (\genblk1.pcpi_mul_mul_2366_47_n_927 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_890 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1413 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48215 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_721 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_828 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_722 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1412 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48217 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_820 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_835 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_425 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1411 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48219 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_788 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_835 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_643 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1410 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48220 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_719 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_835 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_727 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1409 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48221 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_577 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_835 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_534 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1436 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48222 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_755 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_835 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_651 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1408 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48223 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_804 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_835 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_693 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1435 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48224 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_529 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_835 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_479 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1407 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48225 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_256 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_835 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_529 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1434 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48226 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_773 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_835 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_790 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1406 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48227 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_605 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_835 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_417 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1405 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48228 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_764 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_835 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_449 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1433 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48229 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_479 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_835 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_503 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1432 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48230 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_665 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_835 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_403 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1431 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48231 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_613 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_835 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_771 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1404 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48232 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_236 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_836 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_297 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1403 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48233 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_344 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_836 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_331 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1402 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48234 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_331 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_836 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_288 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1401 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48235 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_329 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_836 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_309 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1400 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48236 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_347 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_836 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_268 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1399 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48237 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_457 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_827 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_262 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1398 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48238 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_501 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_829 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_732 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1397 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48239 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_249 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_832 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_807 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1396 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48240 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_646 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_828 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_438 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1395 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48241 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_354 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_829 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_630 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1394 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48242 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_757 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_831 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_710 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1393 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48243 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_421 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_833 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_628 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1392 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48244 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_765 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_831 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_620 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1391 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48245 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_749 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_830 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_263 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1390 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48246 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_580 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_834 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_681 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1389 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48247 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_729 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_825 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_420 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1388 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48248 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_363 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_829 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_714 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1387 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48249 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_674 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_831 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_447 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1386 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48250 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_785 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_828 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_623 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1385 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48251 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_807 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_832 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_609 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1384 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48252 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_629 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_830 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_812 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1383 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48253 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_726 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_834 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_774 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1382 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48254 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_407 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_825 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_428 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1381 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48255 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_447 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_831 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_364 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1380 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48257 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_265 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_824 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_524 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1379 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48258 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_397 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_833 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_742 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1378 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48259 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_766 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_825 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_407 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1377 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48260 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_612 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_831 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_640 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1376 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48261 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_618 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_825 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_655 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1375 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48262 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_388 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_826 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_367 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1374 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48263 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_703 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_831 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_435 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1373 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48264 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_387 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_834 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_813 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1372 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48265 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_779 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_834 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_738 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1371 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48266 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_616 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_825 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_366 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1370 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48267 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_738 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_834 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_580 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1369 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48268 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_692 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_833 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_720 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1368 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48269 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_438 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_828 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_709 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1367 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48270 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_602 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_824 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_723 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1366 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48271 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_600 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_831 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_703 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1365 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48272 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_376 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_825 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_667 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1364 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48273 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_685 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_834 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_779 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1363 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48274 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_734 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_830 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_629 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1362 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48275 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_578 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_830 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_769 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1361 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48276 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_753 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_829 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_772 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1360 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48277 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_671 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_829 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_718 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1359 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48278 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_267 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_831 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_715 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1358 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48279 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_244 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_824 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_679 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1357 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48280 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_489 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_827 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_378 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1356 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48281 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_483 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_831 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_799 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1355 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48282 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_667 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_825 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_616 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1354 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48283 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_760 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_833 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_758 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1353 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48284 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_379 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_832 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_266 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1352 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48285 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_624 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_833 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_585 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1351 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48286 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_382 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_828 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_473 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1350 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48287 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_778 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_828 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_721 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1349 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48288 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_245 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_823 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_731 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1348 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48289 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_450 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_829 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_671 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1347 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48290 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_531 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_832 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_446 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1346 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48291 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_664 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_830 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_743 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1345 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48292 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_634 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_834 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_685 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1344 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48293 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_636 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_833 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_686 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1343 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48294 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_391 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_830 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_801 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1342 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48295 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_663 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_831 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_811 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1341 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48296 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_502 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_825 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_376 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1340 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48297 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_784 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_833 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_636 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1339 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48298 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_617 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_830 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_734 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1338 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48299 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_621 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_830 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_776 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1337 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48300 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_673 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_834 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_726 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1336 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48301 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_425 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_835 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_445 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1335 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48302 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_464 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_831 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_483 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1334 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48303 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_257 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_823 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_638 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1333 ));
  NOR2BX1 \genblk1.pcpi_mul_mul_2366_47_g48304 (.AN
       (\genblk1.pcpi_mul_mul_2366_47_n_928 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_886 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1332 ));
  NOR2BX1 \genblk1.pcpi_mul_mul_2366_47_g48305 (.AN
       (\genblk1.pcpi_mul_mul_2366_47_n_929 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_889 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1331 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48306 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_504 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_825 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_783 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1330 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48307 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_452 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_822 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_713 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1329 ));
  NOR2BX1 \genblk1.pcpi_mul_mul_2366_47_g48308 (.AN
       (\genblk1.pcpi_mul_mul_2366_47_n_918 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_885 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1328 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48309 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_513 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_824 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_414 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1327 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48310 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_731 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_823 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_257 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1326 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48311 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_607 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_826 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_652 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1325 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48312 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_727 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_835 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_613 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1324 ));
  NOR2BX1 \genblk1.pcpi_mul_mul_2366_47_g48313 (.AN
       (\genblk1.pcpi_mul_mul_2366_47_n_924 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_887 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1323 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48314 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_737 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_826 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_649 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1322 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48315 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_583 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_826 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_632 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1321 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48316 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_716 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_835 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_518 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1320 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48317 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_676 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_835 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_719 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1319 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48318 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_364 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_831 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_612 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1318 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48319 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_534 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_835 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_676 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1317 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48320 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_786 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_824 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_756 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1316 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48321 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_751 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_827 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_356 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1315 ));
  NOR2BX1 \genblk1.pcpi_mul_mul_2366_47_g48322 (.AN
       (\genblk1.pcpi_mul_mul_2366_47_n_925 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_882 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1314 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48323 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_769 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_830 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_492 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1313 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48324 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_448 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_830 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_582 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1312 ));
  NOR2BX1 \genblk1.pcpi_mul_mul_2366_47_g48325 (.AN
       (\genblk1.pcpi_mul_mul_2366_47_n_930 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_884 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1311 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48326 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_377 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_834 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_468 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1310 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48327 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_693 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_835 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_577 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1309 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48329 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_768 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_823 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_658 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1308 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48330 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_409 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_833 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_494 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1307 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48331 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_426 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_824 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_265 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1306 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48332 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_699 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_826 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_740 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1305 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48333 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_503 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_835 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_804 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1304 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48334 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_416 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_828 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_759 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1303 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48335 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_741 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_826 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_437 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1302 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48336 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_714 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_829 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_666 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1301 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48337 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_440 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_829 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_800 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1300 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48338 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_518 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_835 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_256 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1299 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48339 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_730 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_822 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_588 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1298 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48340 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_728 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_822 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_791 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1297 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48341 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_650 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_832 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_478 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1296 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48343 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_735 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_829 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_501 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1295 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48344 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_724 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_822 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_452 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1294 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48345 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_625 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_835 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_716 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1293 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48346 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_417 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_835 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_625 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1292 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48347 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_608 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_830 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_639 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1291 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48348 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_414 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_824 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_707 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1290 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48350 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_482 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_827 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_751 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1289 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48351 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_772 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_829 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_363 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1288 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48352 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_771 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_835 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_773 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1287 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48353 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_718 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_829 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_735 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1286 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48354 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_521 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_832 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_650 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1285 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48355 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_651 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_835 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_605 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1284 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48357 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_357 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_835 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_755 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1283 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48358 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_460 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_824 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_474 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1282 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48359 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_262 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_827 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_471 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1281 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48360 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_449 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_835 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_357 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1280 ));
  NOR2BX1 \genblk1.pcpi_mul_mul_2366_47_g48361 (.AN
       (\genblk1.pcpi_mul_mul_2366_47_n_926 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_888 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1279 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48362 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_532 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_822 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_724 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1278 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48363 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_705 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_824 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_513 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1277 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48364 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_647 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_827 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_744 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1276 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48365 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_702 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_826 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_583 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1275 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48366 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_706 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_823 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_490 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1274 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48367 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_643 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_835 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_820 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1273 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48369 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_260 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_826 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_699 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1272 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48370 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_700 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_833 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_515 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1271 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48371 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_403 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_835 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_764 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1270 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48372 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_596 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_824 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_697 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1269 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48373 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_744 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_827 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_712 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1268 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48376 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_537 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_827 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_704 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1267 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48377 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_445 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_835 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_665 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1266 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48378 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_362 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_825 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_766 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1265 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48379 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_395 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_822 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_532 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1264 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48380 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_308 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_836 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_296 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1263 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48381 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_690 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_830 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_586 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1262 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48382 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_343 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_836 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_348 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1261 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48383 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_688 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_823 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_706 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1260 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48384 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_296 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_836 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_300 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1259 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48385 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_686 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_833 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_700 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1258 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48387 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_626 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_827 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_647 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1257 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48388 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_770 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_825 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_255 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1256 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48389 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_278 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_836 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_308 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1255 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48390 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_683 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_827 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_482 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1254 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48391 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_743 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_830 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_608 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1253 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48392 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_323 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_836 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_330 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1252 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48393 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_283 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_836 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_347 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1251 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48394 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_288 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_836 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_329 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1250 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48395 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_678 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_826 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_675 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1249 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48396 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_679 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_824 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_426 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1248 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48397 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_446 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_832 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_521 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1247 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48398 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_628 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_833 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_397 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1246 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48399 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_295 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_836 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_283 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1245 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48400 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_660 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_824 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_705 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1244 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48401 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_309 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_836 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_272 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1243 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48402 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_669 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_826 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_260 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1242 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48405 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_639 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_830 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_448 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1241 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48406 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_477 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_824 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_592 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1240 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48407 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_655 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_825 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_362 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1239 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48408 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_302 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_836 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_278 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1238 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48409 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_304 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_836 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_323 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1237 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48410 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_632 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_826 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_388 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1236 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48411 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_348 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_836 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_302 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1235 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48412 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_495 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_824 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_477 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1234 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48413 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_661 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_828 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_809 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1233 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48414 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_307 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_836 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_789 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1232 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48415 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_748 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_832 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_375 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1231 ));
  NOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48416 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_819 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_891 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1430 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48417 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_310 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_836 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_295 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1230 ));
  NOR2BX1 \genblk1.pcpi_mul_mul_2366_47_g48418 (.AN
       (\genblk1.pcpi_mul_mul_2366_47_n_922 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_883 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1229 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48419 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_275 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_836 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_304 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1228 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48420 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_781 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_828 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_646 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1227 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48421 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_711 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_822 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_395 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1226 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48422 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_648 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_824 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_596 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1225 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48423 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_687 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_826 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_678 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1224 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48424 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_312 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_836 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_343 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1223 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48425 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_630 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_829 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_753 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1222 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48426 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_322 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_836 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_310 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1221 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48427 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_776 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_830 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_690 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1220 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48428 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_645 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_827 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_683 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1219 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48429 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_471 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_827 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_537 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1218 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48430 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_641 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_834 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_673 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1217 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48431 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_470 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_834 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_691 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1216 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48432 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_355 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_826 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_669 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1215 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48433 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_708 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_823 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_688 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1214 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48434 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_332 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_836 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_275 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1213 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48435 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_330 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_836 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_344 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1212 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48436 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_384 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_827 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_626 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1211 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48437 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_811 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_831 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_600 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1210 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48438 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_635 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_824 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_495 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1209 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48439 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_300 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_836 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_322 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1208 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48440 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_297 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_836 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_333 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1207 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48441 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_386 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_828 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_778 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1206 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48442 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_631 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_827 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_384 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1205 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48443 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_333 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_836 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_315 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1204 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48444 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_311 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_836 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_312 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1203 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48445 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_237 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_826 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_355 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1202 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48446 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_486 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_823 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_708 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1201 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48447 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_627 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_826 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_702 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1200 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48448 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_315 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_836 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_311 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1199 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48449 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_622 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_824 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_460 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1198 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48451 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_599 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_832 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_531 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1197 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48452 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_689 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_822 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_711 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1196 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48453 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_268 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_836 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_332 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1195 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48454 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_476 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_824 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_660 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1194 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48455 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_427 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_822 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_728 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1193 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48456 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_292 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_836 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_307 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1192 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48457 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_272 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_836 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_292 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1428 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48458 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_499 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_828 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_762 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1426 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48459 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_698 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_826 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_396 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1424 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48460 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_677 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_827 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_489 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1422 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48461 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_367 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_826 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_741 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1420 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48462 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_715 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_831 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_464 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1418 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48463 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_412 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_822 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_427 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1416 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_g48464 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1189 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1190 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_g48465 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1187 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1188 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_g48466 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1185 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1186 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_g48467 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1183 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1184 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_g48468 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1181 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1182 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_g48469 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1179 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1180 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_g48470 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_1177 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1178 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48471 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_441 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_832 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_606 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1191 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48472 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_242 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_830 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_576 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1176 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48473 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_816 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_825 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_770 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1175 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48474 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_638 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_823 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_668 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1174 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48475 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_390 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_833 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_692 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1173 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48476 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_246 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_828 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_506 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1172 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48477 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_437 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_826 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_694 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1171 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48478 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_424 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_833 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_409 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1170 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48479 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_408 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_832 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_748 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1169 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48480 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_767 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_828 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_781 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1168 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48481 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_253 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_833 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_657 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1167 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48482 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_496 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_833 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_684 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1166 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48483 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_398 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_832 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_797 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1165 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48484 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_523 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_834 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_590 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1164 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48485 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_405 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_822 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_505 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1163 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48486 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_589 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_833 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_784 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1162 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48487 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_413 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_833 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_624 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1161 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48488 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_710 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_831 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_352 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1160 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48489 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_266 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_832 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_408 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1159 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48490 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_587 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_829 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_584 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1158 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48491 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_358 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_831 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_466 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1157 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48492 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_681 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_834 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_603 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1156 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48493 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_439 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_831 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_458 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1155 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48494 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_582 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_830 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_682 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1154 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48495 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_515 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_833 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_717 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1153 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48496 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_239 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_827 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_254 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1152 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48497 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_774 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_834 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_805 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1151 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48498 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_604 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_830 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_662 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1150 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48499 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_389 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_822 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_680 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1149 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48500 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_680 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_822 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_368 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1148 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48501 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_492 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_830 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_604 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1147 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48502 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_240 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_829 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_453 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1146 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48503 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_238 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_825 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_611 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1145 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48504 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_620 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_831 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_358 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1144 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48505 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_780 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_825 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_777 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1143 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48506 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_453 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_829 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_431 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1142 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48507 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_349 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_834 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_641 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1141 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48508 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_691 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_834 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_614 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1140 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48509 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_468 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_834 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_423 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1139 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48510 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_241 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_834 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_517 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1138 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48511 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_623 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_828 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_696 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1137 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48512 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_243 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_822 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_405 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1136 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48513 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_732 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_829 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_353 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1135 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48514 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_261 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_833 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_421 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1134 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48515 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_670 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_830 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_593 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1133 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48516 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_579 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_825 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_504 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1132 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48517 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_436 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_825 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_488 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1131 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48518 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_586 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_830 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_578 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1130 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48519 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_404 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_823 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_653 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1129 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48520 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_666 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_829 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_491 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1128 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48521 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_739 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_831 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_581 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1127 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48522 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_759 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_828 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_402 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1126 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48523 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_465 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_831 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_637 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1125 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48524 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_510 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_829 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_761 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1124 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48525 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_393 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_829 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_633 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1123 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48526 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_662 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_830 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_392 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1122 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48527 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_371 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_832 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_451 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1121 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48528 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_351 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_830 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_670 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1120 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48529 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_508 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_833 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_390 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1119 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48530 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_758 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_833 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_411 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1118 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48531 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_394 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_825 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_594 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1117 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48532 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_506 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_828 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_806 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1116 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48533 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_598 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_825 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_436 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1115 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48534 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_722 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_828 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_785 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1114 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48535 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_512 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_832 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_818 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1113 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48536 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_350 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_832 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_463 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1112 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48537 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_498 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_828 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_499 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1111 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48538 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_682 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_830 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_672 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1110 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48539 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_812 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_830 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_749 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1109 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48540 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_252 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_831 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_739 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1108 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48541 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_469 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_829 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_775 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1107 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48542 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_810 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_822 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_359 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1106 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48543 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_672 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_830 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_617 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1105 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48544 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_777 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_825 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_514 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1104 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48545 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_696 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_828 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_516 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1103 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48546 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_383 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_825 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_502 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1102 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48547 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_640 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_831 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_642 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1101 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48548 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_353 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_829 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_393 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1100 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48549 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_514 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_825 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_816 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1099 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48550 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_754 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_831 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_465 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1098 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48551 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_783 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_825 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_598 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1097 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48552 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_516 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_828 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_507 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1096 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48553 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_752 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_829 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_520 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1095 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48554 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_597 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_832 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_599 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1094 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48555 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_519 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_834 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_349 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1093 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48556 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_511 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_830 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_351 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1092 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48557 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_422 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_825 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_383 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1091 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48558 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_484 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_828 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_695 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1090 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48559 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_633 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_829 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_354 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1089 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48560 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_359 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_822 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_763 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1088 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48561 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_454 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_832 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_372 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1087 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48562 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_411 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_833 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_261 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1086 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48563 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_576 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_830 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_511 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1085 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48564 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_590 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_834 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_470 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1084 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48565 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_642 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_831 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_526 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1083 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48566 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_787 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_823 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_406 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1082 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48567 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_497 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_833 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_413 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1081 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48568 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_381 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_827 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_374 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1080 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48569 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_392 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_830 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_745 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1079 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48570 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_481 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_827 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_677 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1078 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48571 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_675 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_826 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_607 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1077 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48572 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_251 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_831 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_439 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1076 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48573 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_701 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_824 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_817 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1075 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48574 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_584 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_829 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_450 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1074 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48575 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_493 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_822 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_475 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1073 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48576 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_365 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_823 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_793 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1072 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48577 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_475 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_822 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_433 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1071 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48578 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_695 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_828 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_591 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1070 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48579 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_592 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_824 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_385 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1069 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48580 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_707 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_824 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_648 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1068 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48581 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_385 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_824 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_786 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1067 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48582 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_372 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_832 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_512 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1066 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48583 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_520 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_829 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_258 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1065 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48584 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_259 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_823 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_787 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1064 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48585 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_524 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_824 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_527 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1063 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48586 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_500 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_829 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_440 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1062 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48587 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_806 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_828 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_484 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1061 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48588 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_526 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_831 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_252 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1060 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48589 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_588 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_822 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_493 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1059 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48590 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_406 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_823 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_410 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1058 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48591 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_697 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_824 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_380 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1057 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48592 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_756 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_824 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_485 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1056 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48593 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_443 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_827 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_481 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1055 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48594 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_775 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_829 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_752 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1054 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48595 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_463 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_832 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_454 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1053 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48596 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_435 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_831 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_765 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1052 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48597 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_750 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_834 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_794 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1051 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48598 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_611 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_825 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_394 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1050 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48599 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_472 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_834 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_523 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1049 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48600 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_533 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_823 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_365 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1048 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48601 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_594 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_825 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_579 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1047 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48602 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_517 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_834 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_377 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1046 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48603 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_535 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_826 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_802 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1045 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48604 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_370 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_827 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_381 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1044 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48605 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_466 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_831 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_754 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1043 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48606 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_709 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_828 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_416 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1042 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48607 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_442 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_832 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_455 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1041 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48608 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_536 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_826 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_595 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1040 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48609 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_509 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_825 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_422 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1039 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48610 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_813 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_834 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_472 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1038 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48611 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_410 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_823 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_429 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1037 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48612 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_254 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_827 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_456 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1036 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48613 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_375 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_832 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_399 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1035 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48614 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_380 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_824 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_622 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1034 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48615 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_462 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_823 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_259 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1033 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48616 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_485 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_824 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_476 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1032 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48617 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_418 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_823 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_462 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1031 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48618 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_725 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_822 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_730 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1030 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48619 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_451 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_832 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_350 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1029 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48620 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_401 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_832 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_442 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1028 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48621 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_528 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_827 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_457 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1027 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48622 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_694 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_826 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_698 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1026 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48623 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_433 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_822 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_530 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1025 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48624 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_415 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_834 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_750 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1024 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48625 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_461 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_824 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_701 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1023 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48626 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_614 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_834 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_736 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1022 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48627 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_258 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_829 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_419 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1021 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48628 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_591 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_828 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_814 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1020 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48629 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_615 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_826 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_737 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1019 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48630 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_430 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_823 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_747 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1018 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48631 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_494 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_833 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_497 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1017 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48632 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_712 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_827 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_487 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1016 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48633 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_601 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_823 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_361 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1015 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48634 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_444 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_822 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_725 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1014 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48635 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_653 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_823 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_418 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1013 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48636 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_809 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_828 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_382 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1012 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48637 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_746 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_834 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_387 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1011 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48638 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_619 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_832 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_371 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1010 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48639 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_263 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_830 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_391 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1009 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48640 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_742 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_833 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_424 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1008 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48641 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_369 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_822 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_444 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1007 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48642 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_455 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_832 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_398 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1006 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48643 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_456 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_827 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_808 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1005 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48644 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_659 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_826 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_733 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1004 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48645 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_423 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_834 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_746 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1003 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48646 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_818 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_832 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_597 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1002 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48647 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_530 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_822 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_480 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1001 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48648 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_814 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_828 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_767 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1000 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48649 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_740 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_826 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_656 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_999 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48650 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_473 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_828 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_795 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_998 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48651 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_654 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_823 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_404 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_997 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48652 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_704 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_827 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_803 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_996 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48653 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_763 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_822 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_412 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_995 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48654 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_434 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_822 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_369 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_994 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48655 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_264 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_832 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_619 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_993 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48656 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_717 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_833 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_400 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_992 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48657 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_419 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_829 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_587 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_991 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48658 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_736 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_834 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_634 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_990 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48659 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_723 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_824 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_796 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_989 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48660 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_459 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_823 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_533 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_988 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48661 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_429 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_823 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_815 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_987 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48662 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_248 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_833 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_589 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_986 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48663 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_782 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_827 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_443 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_985 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48664 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_368 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_822 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_434 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_984 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48665 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_762 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_828 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_386 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_983 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48666 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_361 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_823 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_654 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_982 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48667 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_402 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_828 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_525 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_981 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48668 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_399 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_832 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_264 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_980 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48669 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_713 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_822 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_373 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_979 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48670 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_745 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_830 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_664 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_978 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48671 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_684 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_833 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_798 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_977 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48672 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_396 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_826 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_535 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_976 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48673 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_428 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_825 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_729 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_975 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48674 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_610 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_826 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_615 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_974 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48675 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_815 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_823 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_486 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_973 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48676 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_467 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_827 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_370 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_972 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48677 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_606 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_832 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_401 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_971 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48678 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_817 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_824 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_635 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_970 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48679 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_637 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_831 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_267 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_969 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48680 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_525 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_828 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_498 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_968 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48681 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_373 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_822 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_810 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_967 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48682 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_747 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_823 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_601 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_966 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48683 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_656 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_826 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_610 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_965 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48684 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_649 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_826 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_687 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_964 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48685 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_432 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_822 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_389 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_963 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48686 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_527 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_824 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_461 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_962 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48687 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_356 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_827 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_782 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_961 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48688 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_733 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_826 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_536 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_960 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48689 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_658 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_823 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_459 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_959 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48690 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_431 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_829 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_510 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_958 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48691 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_400 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_833 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_760 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_957 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48692 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_652 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_826 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_659 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_956 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48693 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_458 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_831 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_757 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_955 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48694 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_505 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_822 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_432 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_954 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48695 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_366 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_825 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_780 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_953 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48696 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_603 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_834 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_360 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_952 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48697 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_374 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_827 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_645 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_951 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48698 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_487 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_827 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_467 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_950 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48699 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_522 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_823 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_430 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_949 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48700 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_490 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_823 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_768 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_948 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48701 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_480 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_822 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_689 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_947 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48702 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_644 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_823 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_522 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_946 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48703 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_488 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_825 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_618 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_945 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48704 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_255 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_825 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_792 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_944 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48705 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_352 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_831 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_674 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_943 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48706 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_761 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_829 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_469 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_942 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48707 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_360 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_834 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_519 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_941 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48708 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_378 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_827 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_528 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_940 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48709 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_581 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_831 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_663 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_939 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48710 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_808 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_827 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_631 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_938 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48711 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_478 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_832 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_441 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_937 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48712 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_507 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_828 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_661 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_936 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48713 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_593 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_830 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_621 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_935 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48714 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_609 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_832 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_379 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_934 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48715 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_595 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_826 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_627 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_933 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48716 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_668 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_823 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_644 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_932 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48717 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_491 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_829 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_500 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1189 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48718 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_585 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_833 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_253 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1187 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48719 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_720 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_833 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_496 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1185 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48720 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_805 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_834 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_415 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1183 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48721 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_657 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_833 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_508 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1181 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48722 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_420 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_825 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_509 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1179 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48723 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_474 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_824 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_602 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1177 ));
  NOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48724 (.A
       (\genblk1.pcpi_mul_rs1 [0]), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_226 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_931 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48725 (.A0
       (\genblk1.pcpi_mul_rs2 [29]), .A1 (n_11757), .B0
       (\genblk1.pcpi_mul_rs2 [30]), .B1 (\genblk1.pcpi_mul_rs1 [0]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_930 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48726 (.A0
       (\genblk1.pcpi_mul_rs2 [11]), .A1 (n_11756), .B0
       (\genblk1.pcpi_mul_rs2 [12]), .B1 (\genblk1.pcpi_mul_rs1 [0]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_196 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_929 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48727 (.A0
       (\genblk1.pcpi_mul_rs2 [15]), .A1 (n_11751), .B0
       (\genblk1.pcpi_mul_rs2 [16]), .B1 (\genblk1.pcpi_mul_rs1 [0]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_194 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_928 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48728 (.A0
       (\genblk1.pcpi_mul_rs2 [1]), .A1 (n_11750), .B0
       (\genblk1.pcpi_mul_rs1 [0]), .B1 (\genblk1.pcpi_mul_rs2 [2]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_165 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_927 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48729 (.A0
       (\genblk1.pcpi_mul_rs2 [27]), .A1 (n_11755), .B0
       (\genblk1.pcpi_mul_rs2 [28]), .B1 (\genblk1.pcpi_mul_rs1 [0]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_197 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_926 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48730 (.A0
       (\genblk1.pcpi_mul_rs2 [13]), .A1 (n_11758), .B0
       (\genblk1.pcpi_mul_rs2 [14]), .B1 (\genblk1.pcpi_mul_rs1 [0]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_166 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_925 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48731 (.A0
       (\genblk1.pcpi_mul_rs2 [3]), .A1 (n_11754), .B0
       (\genblk1.pcpi_mul_rs2 [4]), .B1 (\genblk1.pcpi_mul_rs1 [0]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_170 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_924 ));
  OAI211X1 \genblk1.pcpi_mul_mul_2366_47_g48732 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_14 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .B0
       (\genblk1.pcpi_mul_rs2 [9]), .C0
       (\genblk1.pcpi_mul_mul_2366_47_n_558 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_923 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48733 (.A0
       (\genblk1.pcpi_mul_rs2 [5]), .A1 (n_11752), .B0
       (\genblk1.pcpi_mul_rs2 [6]), .B1 (\genblk1.pcpi_mul_rs1 [0]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_167 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_922 ));
  OAI211X1 \genblk1.pcpi_mul_mul_2366_47_g48734 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_16 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .B0
       (\genblk1.pcpi_mul_rs2 [25]), .C0
       (\genblk1.pcpi_mul_mul_2366_47_n_539 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_921 ));
  OAI211X1 \genblk1.pcpi_mul_mul_2366_47_g48735 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_22 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .B0
       (\genblk1.pcpi_mul_rs2 [27]), .C0
       (\genblk1.pcpi_mul_mul_2366_47_n_557 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_920 ));
  OAI211X1 \genblk1.pcpi_mul_mul_2366_47_g48736 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_18 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .B0
       (\genblk1.pcpi_mul_rs2 [23]), .C0
       (\genblk1.pcpi_mul_mul_2366_47_n_556 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_919 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48737 (.A0
       (\genblk1.pcpi_mul_rs2 [17]), .A1 (n_11753), .B0
       (\genblk1.pcpi_mul_rs2 [18]), .B1 (\genblk1.pcpi_mul_rs1 [0]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_164 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_918 ));
  OAI211X1 \genblk1.pcpi_mul_mul_2366_47_g48738 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_20 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .B0
       (\genblk1.pcpi_mul_rs2 [21]), .C0
       (\genblk1.pcpi_mul_mul_2366_47_n_555 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_917 ));
  OAI211X1 \genblk1.pcpi_mul_mul_2366_47_g48739 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_24 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .B0
       (\genblk1.pcpi_mul_rs2 [11]), .C0
       (\genblk1.pcpi_mul_mul_2366_47_n_554 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_916 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48740 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_172 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_81 ), .B0
       (\genblk1.pcpi_mul_rs2 [32]), .B1 (\genblk1.pcpi_mul_rs1 [1]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_137 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_915 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48741 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_172 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_71 ), .B0
       (\genblk1.pcpi_mul_rs2 [32]), .B1 (\genblk1.pcpi_mul_rs1 [4]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_137 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_914 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48742 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_172 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_75 ), .B0
       (\genblk1.pcpi_mul_rs2 [32]), .B1 (\genblk1.pcpi_mul_rs1 [9]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_137 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_913 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48743 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_73 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_172 ), .B0
       (\genblk1.pcpi_mul_rs1 [19]), .B1 (\genblk1.pcpi_mul_rs2 [32]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_137 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_912 ));
  NOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48744 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_137 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_911 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48745 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_53 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_172 ), .B0
       (\genblk1.pcpi_mul_rs1 [25]), .B1 (\genblk1.pcpi_mul_rs2 [32]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_137 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_910 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48746 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_67 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_172 ), .B0
       (\genblk1.pcpi_mul_rs1 [21]), .B1 (\genblk1.pcpi_mul_rs2 [32]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_137 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_909 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48747 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_172 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_91 ), .B0
       (\genblk1.pcpi_mul_rs2 [32]), .B1 (\genblk1.pcpi_mul_rs1 [7]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_137 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_908 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48748 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_99 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_172 ), .B0
       (\genblk1.pcpi_mul_rs1 [24]), .B1 (\genblk1.pcpi_mul_rs2 [32]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_137 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_907 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48749 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_172 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_57 ), .B0
       (\genblk1.pcpi_mul_rs2 [32]), .B1 (\genblk1.pcpi_mul_rs1 [2]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_137 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_906 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48750 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_172 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_39 ), .B0
       (\genblk1.pcpi_mul_rs2 [32]), .B1 (\genblk1.pcpi_mul_rs1 [14]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_137 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_905 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48751 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_87 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_172 ), .B0
       (\genblk1.pcpi_mul_rs1 [20]), .B1 (\genblk1.pcpi_mul_rs2 [32]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_137 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_904 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48752 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_172 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_69 ), .B0
       (\genblk1.pcpi_mul_rs2 [32]), .B1 (\genblk1.pcpi_mul_rs1 [10]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_137 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_903 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48753 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_172 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_51 ), .B0
       (\genblk1.pcpi_mul_rs2 [32]), .B1 (\genblk1.pcpi_mul_rs1 [11]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_137 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_902 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48754 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_172 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_83 ), .B0
       (\genblk1.pcpi_mul_rs2 [32]), .B1 (\genblk1.pcpi_mul_rs1 [17]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_137 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_901 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48755 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_172 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_59 ), .B0
       (\genblk1.pcpi_mul_rs2 [32]), .B1 (\genblk1.pcpi_mul_rs1 [6]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_137 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_900 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48756 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_172 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_97 ), .B0
       (\genblk1.pcpi_mul_rs2 [32]), .B1 (\genblk1.pcpi_mul_rs1 [15]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_137 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_899 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48757 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_49 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_172 ), .B0
       (\genblk1.pcpi_mul_rs1 [23]), .B1 (\genblk1.pcpi_mul_rs2 [32]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_137 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_898 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48758 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_61 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_172 ), .B0
       (\genblk1.pcpi_mul_rs1 [29]), .B1 (\genblk1.pcpi_mul_rs2 [32]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_137 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_897 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48759 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_172 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_47 ), .B0
       (\genblk1.pcpi_mul_rs2 [32]), .B1 (\genblk1.pcpi_mul_rs1 [5]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_137 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_896 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48760 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_77 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_172 ), .B0
       (\genblk1.pcpi_mul_rs1 [27]), .B1 (\genblk1.pcpi_mul_rs2 [32]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_137 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_895 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48761 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_79 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_172 ), .B0
       (\genblk1.pcpi_mul_rs1 [18]), .B1 (\genblk1.pcpi_mul_rs2 [32]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_137 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_894 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48762 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_172 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_45 ), .B0
       (\genblk1.pcpi_mul_rs2 [32]), .B1 (\genblk1.pcpi_mul_rs1 [12]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_137 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_893 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48763 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_172 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_93 ), .B0
       (\genblk1.pcpi_mul_rs2 [32]), .B1 (\genblk1.pcpi_mul_rs1 [3]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_137 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_892 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48764 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_223 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_250 ), .B0
       (\genblk1.pcpi_mul_rs2 [0]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_279 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_891 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48765 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_224 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_280 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_35 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_327 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_880 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48766 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_43 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_172 ), .B0
       (\genblk1.pcpi_mul_rs1 [31]), .B1 (\genblk1.pcpi_mul_rs2 [32]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_137 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_879 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48767 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_223 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_328 ), .B0
       (\genblk1.pcpi_mul_rs2 [0]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_334 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_890 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48768 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_223 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_271 ), .B0
       (\genblk1.pcpi_mul_rs2 [0]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_305 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_889 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48769 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_223 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_294 ), .B0
       (\genblk1.pcpi_mul_rs2 [0]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_276 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_888 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48770 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_223 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_314 ), .B0
       (\genblk1.pcpi_mul_rs2 [0]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_338 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_887 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48771 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_223 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_274 ), .B0
       (\genblk1.pcpi_mul_rs2 [0]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_298 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_886 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48772 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_223 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_342 ), .B0
       (\genblk1.pcpi_mul_rs2 [0]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_318 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_885 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48773 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_223 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_289 ), .B0
       (\genblk1.pcpi_mul_rs2 [0]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_324 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_884 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48774 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_223 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_346 ), .B0
       (\genblk1.pcpi_mul_rs2 [0]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_320 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_883 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48775 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_223 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_287 ), .B0
       (\genblk1.pcpi_mul_rs2 [0]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_281 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_882 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48776 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_172 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_41 ), .B0
       (\genblk1.pcpi_mul_rs2 [32]), .B1 (\genblk1.pcpi_mul_rs1 [13]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_137 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_878 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48777 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_224 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_317 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_35 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_270 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_877 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48778 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_224 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_335 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_35 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_313 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_876 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48779 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_224 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_336 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_35 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_285 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_875 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48780 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_224 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_340 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_35 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_336 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_874 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48781 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_55 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_172 ), .B0
       (\genblk1.pcpi_mul_rs1 [26]), .B1 (\genblk1.pcpi_mul_rs2 [32]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_137 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_873 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48782 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_224 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_277 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_35 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_290 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_872 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48783 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_224 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_325 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_35 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_538 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_871 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48784 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_224 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_306 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_35 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_286 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_870 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48785 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_95 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_172 ), .B0
       (\genblk1.pcpi_mul_rs1 [22]), .B1 (\genblk1.pcpi_mul_rs2 [32]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_137 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_869 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48786 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_224 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_326 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_35 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_293 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_868 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48787 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_224 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_321 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_35 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_340 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_867 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48788 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_224 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_337 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_35 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_326 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_866 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48789 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_224 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_291 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_35 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_316 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_865 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48790 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_224 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_284 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_35 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_291 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_864 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48791 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_224 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_269 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_35 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_284 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_863 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48792 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_89 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_172 ), .B0
       (\genblk1.pcpi_mul_rs2 [32]), .B1 (\genblk1.pcpi_mul_rs1 [16]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_137 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_862 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48793 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_224 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_303 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_35 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_301 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_861 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48794 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_172 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_85 ), .B0
       (\genblk1.pcpi_mul_rs2 [32]), .B1 (\genblk1.pcpi_mul_rs1 [8]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_137 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_860 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48795 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_224 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_319 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_35 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_303 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_859 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48796 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_224 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_339 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_35 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_345 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_858 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48797 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_224 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_316 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_35 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_337 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_857 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48798 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_224 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_282 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_35 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_273 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_856 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48799 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_224 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_299 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_35 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_341 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_855 ));
  AOI221X1 \genblk1.pcpi_mul_mul_2366_47_g48800 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_65 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_172 ), .B0
       (\genblk1.pcpi_mul_rs1 [28]), .B1 (\genblk1.pcpi_mul_rs2 [32]),
       .C0 (\genblk1.pcpi_mul_mul_2366_47_n_137 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_854 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48801 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_224 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_285 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_35 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_317 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_853 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48802 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_224 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_301 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_35 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_269 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_852 ));
  OAI221X1 \genblk1.pcpi_mul_mul_2366_47_g48803 (.A0
       (\genblk1.pcpi_mul_rs1 [30]), .A1 (\genblk1.pcpi_mul_rs2 [32]),
       .B0 (\genblk1.pcpi_mul_mul_2366_47_n_63 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_172 ), .C0
       (\genblk1.pcpi_mul_mul_2366_47_n_162 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_881 ));
  NOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48805 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_851 ));
  NOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48806 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_850 ));
  NOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48807 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_849 ));
  NOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48808 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_848 ));
  NOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48809 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_847 ));
  NOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48810 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_846 ));
  NOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48811 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_845 ));
  NOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48812 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_844 ));
  NOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48813 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_843 ));
  NOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48814 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_842 ));
  NOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48815 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_841 ));
  NOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48816 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_840 ));
  NOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48817 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_839 ));
  NOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48818 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_838 ));
  NOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48819 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_837 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48820 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_228 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_227 ), .B0
       (\genblk1.pcpi_mul_rs2 [0]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_223 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_821 ));
  OR2X2 \genblk1.pcpi_mul_mul_2366_47_g48821 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_553 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_156 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_836 ));
  OR2X2 \genblk1.pcpi_mul_mul_2366_47_g48822 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_547 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_148 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_835 ));
  OR2X2 \genblk1.pcpi_mul_mul_2366_47_g48823 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_540 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_147 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_834 ));
  OR2X2 \genblk1.pcpi_mul_mul_2366_47_g48824 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_552 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_157 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_833 ));
  OR2X2 \genblk1.pcpi_mul_mul_2366_47_g48825 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_551 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_155 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_832 ));
  OR2X2 \genblk1.pcpi_mul_mul_2366_47_g48826 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_542 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_160 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_831 ));
  OR2X2 \genblk1.pcpi_mul_mul_2366_47_g48827 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_548 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_152 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_830 ));
  OR2X2 \genblk1.pcpi_mul_mul_2366_47_g48828 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_546 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_151 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_829 ));
  OR2X2 \genblk1.pcpi_mul_mul_2366_47_g48829 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_544 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_154 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_828 ));
  OR2X2 \genblk1.pcpi_mul_mul_2366_47_g48830 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_543 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_150 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_827 ));
  OR2X2 \genblk1.pcpi_mul_mul_2366_47_g48831 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_545 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_161 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_826 ));
  OR2X2 \genblk1.pcpi_mul_mul_2366_47_g48832 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_559 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_158 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_825 ));
  OR2X2 \genblk1.pcpi_mul_mul_2366_47_g48833 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_541 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_149 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_824 ));
  OR2X2 \genblk1.pcpi_mul_mul_2366_47_g48834 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_549 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_159 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_823 ));
  OR2X2 \genblk1.pcpi_mul_mul_2366_47_g48835 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_550 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_153 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_822 ));
  XNOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48865 (.A
       (\genblk1.pcpi_mul_rs2 [16]), .B (\genblk1.pcpi_mul_rs2 [17]),
       .Y (\genblk1.pcpi_mul_mul_2366_47_n_559 ));
  OAI2BB1X1 \genblk1.pcpi_mul_mul_2366_47_g48866 (.A0N
       (\genblk1.pcpi_mul_mul_2366_47_n_14 ), .A1N
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .B0
       (\genblk1.pcpi_mul_rs2 [7]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_558 ));
  OAI2BB1X1 \genblk1.pcpi_mul_mul_2366_47_g48867 (.A0N
       (\genblk1.pcpi_mul_mul_2366_47_n_22 ), .A1N
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .B0
       (\genblk1.pcpi_mul_rs2 [25]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_557 ));
  OAI2BB1X1 \genblk1.pcpi_mul_mul_2366_47_g48868 (.A0N
       (\genblk1.pcpi_mul_mul_2366_47_n_18 ), .A1N
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .B0
       (\genblk1.pcpi_mul_rs2 [21]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_556 ));
  OAI2BB1X1 \genblk1.pcpi_mul_mul_2366_47_g48869 (.A0N
       (\genblk1.pcpi_mul_mul_2366_47_n_20 ), .A1N
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .B0
       (\genblk1.pcpi_mul_rs2 [19]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_555 ));
  OAI2BB1X1 \genblk1.pcpi_mul_mul_2366_47_g48870 (.A0N
       (\genblk1.pcpi_mul_mul_2366_47_n_24 ), .A1N
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .B0
       (\genblk1.pcpi_mul_rs2 [9]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_554 ));
  XNOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48871 (.A
       (\genblk1.pcpi_mul_rs2 [31]), .B (\genblk1.pcpi_mul_rs2 [30]),
       .Y (\genblk1.pcpi_mul_mul_2366_47_n_553 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48872 (.A0
       (\genblk1.pcpi_mul_rs2 [25]), .A1 (\genblk1.pcpi_mul_rs2 [24]),
       .B0 (\genblk1.pcpi_mul_mul_2366_47_n_198 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_16 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_552 ));
  XNOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48873 (.A
       (\genblk1.pcpi_mul_rs2 [6]), .B (\genblk1.pcpi_mul_rs2 [7]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_551 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48874 (.A0
       (\genblk1.pcpi_mul_rs2 [9]), .A1 (\genblk1.pcpi_mul_rs2 [8]),
       .B0 (\genblk1.pcpi_mul_mul_2366_47_n_163 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_14 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_550 ));
  XNOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48875 (.A
       (\genblk1.pcpi_mul_rs2 [4]), .B (\genblk1.pcpi_mul_rs2 [5]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_549 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48876 (.A0
       (\genblk1.pcpi_mul_rs2 [21]), .A1 (\genblk1.pcpi_mul_rs2 [20]),
       .B0 (\genblk1.pcpi_mul_mul_2366_47_n_195 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_20 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_548 ));
  XNOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48877 (.A
       (\genblk1.pcpi_mul_rs2 [2]), .B (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_547 ));
  XNOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48878 (.A
       (\genblk1.pcpi_mul_rs2 [15]), .B (\genblk1.pcpi_mul_rs2 [14]),
       .Y (\genblk1.pcpi_mul_mul_2366_47_n_546 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48879 (.A0
       (\genblk1.pcpi_mul_rs2 [27]), .A1 (\genblk1.pcpi_mul_rs2 [26]),
       .B0 (\genblk1.pcpi_mul_mul_2366_47_n_193 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_22 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_545 ));
  XNOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48880 (.A
       (\genblk1.pcpi_mul_rs2 [18]), .B (\genblk1.pcpi_mul_rs2 [19]),
       .Y (\genblk1.pcpi_mul_mul_2366_47_n_544 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48881 (.A0
       (\genblk1.pcpi_mul_rs2 [22]), .A1 (\genblk1.pcpi_mul_rs2 [23]),
       .B0 (\genblk1.pcpi_mul_mul_2366_47_n_18 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_543 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g48882 (.A0
       (\genblk1.pcpi_mul_rs2 [10]), .A1 (\genblk1.pcpi_mul_rs2 [11]),
       .B0 (\genblk1.pcpi_mul_mul_2366_47_n_24 ), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_542 ));
  XNOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48883 (.A
       (\genblk1.pcpi_mul_rs2 [28]), .B (\genblk1.pcpi_mul_rs2 [29]),
       .Y (\genblk1.pcpi_mul_mul_2366_47_n_541 ));
  XNOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48884 (.A
       (\genblk1.pcpi_mul_rs2 [13]), .B (\genblk1.pcpi_mul_rs2 [12]),
       .Y (\genblk1.pcpi_mul_mul_2366_47_n_540 ));
  OAI2BB1X1 \genblk1.pcpi_mul_mul_2366_47_g48885 (.A0N
       (\genblk1.pcpi_mul_mul_2366_47_n_16 ), .A1N
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .B0
       (\genblk1.pcpi_mul_rs2 [23]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_539 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48886 (.A0
       (\genblk1.pcpi_mul_rs1 [3]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_165 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_93 ), .B1
       (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_820 ));
  NAND2BX1 \genblk1.pcpi_mul_mul_2366_47_g48887 (.AN
       (\genblk1.pcpi_mul_n_91 ), .B (\genblk1.pcpi_mul_rs2 [1]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_819 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48888 (.A0
       (\genblk1.pcpi_mul_rs1 [18]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_167 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_79 ), .B1
       (\genblk1.pcpi_mul_rs2 [7]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_818 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48889 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_197 ), .A1
       (\genblk1.pcpi_mul_rs1 [8]), .B0 (\genblk1.pcpi_mul_rs2 [29]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_85 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_817 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48890 (.A0
       (\genblk1.pcpi_mul_rs1 [29]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_194 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_61 ), .B1
       (\genblk1.pcpi_mul_rs2 [17]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_816 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48891 (.A0
       (\genblk1.pcpi_mul_rs1 [21]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_170 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_67 ), .B1
       (\genblk1.pcpi_mul_rs2 [5]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_815 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48892 (.A0
       (\genblk1.pcpi_mul_rs1 [6]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_164 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_59 ), .B1
       (\genblk1.pcpi_mul_rs2 [19]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_814 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48893 (.A0
       (\genblk1.pcpi_mul_rs1 [7]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_196 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_91 ), .B1
       (\genblk1.pcpi_mul_rs2 [13]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_813 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48894 (.A0
       (\genblk1.pcpi_mul_rs1 [28]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_195 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_65 ), .B1
       (\genblk1.pcpi_mul_rs2 [21]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_812 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48895 (.A0
       (\genblk1.pcpi_mul_rs1 [17]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_83 ), .B1
       (\genblk1.pcpi_mul_rs2 [11]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_811 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48896 (.A0
       (\genblk1.pcpi_mul_rs1 [26]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_163 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_55 ), .B1
       (\genblk1.pcpi_mul_rs2 [9]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_810 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48897 (.A0
       (\genblk1.pcpi_mul_rs1 [29]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_164 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_61 ), .B1
       (\genblk1.pcpi_mul_rs2 [19]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_809 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48898 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ), .A1
       (\genblk1.pcpi_mul_rs1 [3]), .B0 (\genblk1.pcpi_mul_rs2 [23]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_93 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_808 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48899 (.A0
       (\genblk1.pcpi_mul_rs1 [1]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_167 ), .B0
       (\genblk1.pcpi_mul_rs2 [7]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_81 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_807 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48900 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_164 ), .A1
       (\genblk1.pcpi_mul_rs1 [2]), .B0 (\genblk1.pcpi_mul_rs2 [19]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_57 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_806 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48901 (.A0
       (\genblk1.pcpi_mul_rs1 [29]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_196 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_61 ), .B1
       (\genblk1.pcpi_mul_rs2 [13]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_805 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48902 (.A0
       (\genblk1.pcpi_mul_rs1 [22]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_165 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_95 ), .B1
       (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_804 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48903 (.A0
       (\genblk1.pcpi_mul_rs1 [32]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_37 ), .B1
       (\genblk1.pcpi_mul_rs2 [23]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_803 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48904 (.A0
       (\genblk1.pcpi_mul_rs1 [32]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_193 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_37 ), .B1
       (\genblk1.pcpi_mul_rs2 [27]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_802 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48905 (.A0
       (\genblk1.pcpi_mul_rs1 [32]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_195 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_37 ), .B1
       (\genblk1.pcpi_mul_rs2 [21]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_801 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48906 (.A0
       (\genblk1.pcpi_mul_rs1 [32]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_166 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_37 ), .B1
       (\genblk1.pcpi_mul_rs2 [15]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_800 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48907 (.A0
       (\genblk1.pcpi_mul_rs1 [32]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_37 ), .B1
       (\genblk1.pcpi_mul_rs2 [11]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_799 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48908 (.A0
       (\genblk1.pcpi_mul_rs1 [32]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_198 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_37 ), .B1
       (\genblk1.pcpi_mul_rs2 [25]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_798 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48909 (.A0
       (\genblk1.pcpi_mul_rs1 [32]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_167 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_37 ), .B1
       (\genblk1.pcpi_mul_rs2 [7]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_797 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48910 (.A0
       (\genblk1.pcpi_mul_rs1 [32]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_197 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_37 ), .B1
       (\genblk1.pcpi_mul_rs2 [29]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_796 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48911 (.A0
       (\genblk1.pcpi_mul_rs1 [32]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_164 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_37 ), .B1
       (\genblk1.pcpi_mul_rs2 [19]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_795 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48912 (.A0
       (\genblk1.pcpi_mul_rs1 [32]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_196 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_37 ), .B1
       (\genblk1.pcpi_mul_rs2 [13]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_794 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48913 (.A0
       (\genblk1.pcpi_mul_rs1 [32]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_170 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_37 ), .B1
       (\genblk1.pcpi_mul_rs2 [5]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_793 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48914 (.A0
       (\genblk1.pcpi_mul_rs1 [32]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_194 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_37 ), .B1
       (\genblk1.pcpi_mul_rs2 [17]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_792 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48915 (.A0
       (\genblk1.pcpi_mul_rs1 [32]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_163 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_37 ), .B1
       (\genblk1.pcpi_mul_rs2 [9]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_791 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48916 (.A0
       (\genblk1.pcpi_mul_rs1 [32]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_165 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_37 ), .B1
       (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_790 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48917 (.A0
       (\genblk1.pcpi_mul_rs1 [32]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_37 ), .B1
       (\genblk1.pcpi_mul_rs2 [31]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_789 ));
  NOR2X1 \genblk1.pcpi_mul_mul_2366_47_g48918 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_228 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_227 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_538 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48919 (.A0
       (\genblk1.pcpi_mul_rs1 [1]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_165 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_81 ), .B1
       (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_788 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48920 (.A0
       (\genblk1.pcpi_mul_rs1 [17]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_170 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_83 ), .B1
       (\genblk1.pcpi_mul_rs2 [5]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_787 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48921 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_197 ), .A1
       (\genblk1.pcpi_mul_rs1 [14]), .B0 (\genblk1.pcpi_mul_rs2 [29]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_39 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_786 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48922 (.A0
       (\genblk1.pcpi_mul_rs1 [23]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_164 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_49 ), .B1
       (\genblk1.pcpi_mul_rs2 [19]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_785 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48923 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_198 ), .A1
       (\genblk1.pcpi_mul_rs1 [2]), .B0 (\genblk1.pcpi_mul_rs2 [25]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_57 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_784 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48924 (.A0
       (\genblk1.pcpi_mul_rs1 [6]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_194 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_59 ), .B1
       (\genblk1.pcpi_mul_rs2 [17]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_783 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48925 (.A0
       (\genblk1.pcpi_mul_rs1 [20]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_87 ), .B1
       (\genblk1.pcpi_mul_rs2 [23]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_782 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48926 (.A0
       (\genblk1.pcpi_mul_rs1 [8]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_164 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_85 ), .B1
       (\genblk1.pcpi_mul_rs2 [19]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_781 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48927 (.A0
       (\genblk1.pcpi_mul_rs1 [26]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_194 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_55 ), .B1
       (\genblk1.pcpi_mul_rs2 [17]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_780 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48928 (.A0
       (\genblk1.pcpi_mul_rs1 [17]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_196 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_83 ), .B1
       (\genblk1.pcpi_mul_rs2 [13]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_779 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48929 (.A0
       (\genblk1.pcpi_mul_rs1 [20]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_164 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_87 ), .B1
       (\genblk1.pcpi_mul_rs2 [19]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_778 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48930 (.A0
       (\genblk1.pcpi_mul_rs1 [27]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_194 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_77 ), .B1
       (\genblk1.pcpi_mul_rs2 [17]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_777 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48931 (.A0
       (\genblk1.pcpi_mul_rs1 [7]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_195 ), .B0
       (\genblk1.pcpi_mul_rs2 [21]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_91 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_776 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48932 (.A0
       (\genblk1.pcpi_mul_rs1 [6]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_166 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_59 ), .B1
       (\genblk1.pcpi_mul_rs2 [15]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_775 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48933 (.A0
       (\genblk1.pcpi_mul_rs1 [28]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_196 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_65 ), .B1
       (\genblk1.pcpi_mul_rs2 [13]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_774 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48934 (.A0
       (\genblk1.pcpi_mul_rs1 [31]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_165 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_43 ), .B1
       (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_773 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48935 (.A0
       (\genblk1.pcpi_mul_rs1 [25]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_166 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_53 ), .B1
       (\genblk1.pcpi_mul_rs2 [15]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_772 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48936 (.A0
       (\genblk1.pcpi_mul_rs1 [30]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_165 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_63 ), .B1
       (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_771 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48937 (.A0
       (\genblk1.pcpi_mul_rs1 [30]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_194 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_63 ), .B1
       (\genblk1.pcpi_mul_rs2 [17]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_770 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48938 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_195 ), .A1
       (\genblk1.pcpi_mul_rs1 [11]), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_51 ), .B1
       (\genblk1.pcpi_mul_rs2 [21]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_769 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48939 (.A0
       (\genblk1.pcpi_mul_rs1 [27]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_170 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_77 ), .B1
       (\genblk1.pcpi_mul_rs2 [5]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_768 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48940 (.A0
       (\genblk1.pcpi_mul_rs1 [7]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_164 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_91 ), .B1
       (\genblk1.pcpi_mul_rs2 [19]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_767 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48941 (.A0
       (\genblk1.pcpi_mul_rs1 [13]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_194 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_41 ), .B1
       (\genblk1.pcpi_mul_rs2 [17]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_766 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48942 (.A0
       (\genblk1.pcpi_mul_rs1 [21]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_67 ), .B1
       (\genblk1.pcpi_mul_rs2 [11]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_765 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48943 (.A0
       (\genblk1.pcpi_mul_rs1 [8]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_165 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_85 ), .B1
       (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_764 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48944 (.A0
       (\genblk1.pcpi_mul_rs1 [28]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_163 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_65 ), .B1
       (\genblk1.pcpi_mul_rs2 [9]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_763 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48945 (.A0
       (\genblk1.pcpi_mul_rs1 [18]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_164 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_79 ), .B1
       (\genblk1.pcpi_mul_rs2 [19]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_762 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48946 (.A0
       (\genblk1.pcpi_mul_rs1 [4]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_166 ), .B0
       (\genblk1.pcpi_mul_rs2 [15]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_71 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_761 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48947 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_198 ), .A1
       (\genblk1.pcpi_mul_rs1 [9]), .B0 (\genblk1.pcpi_mul_rs2 [25]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_75 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_760 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48948 (.A0
       (\genblk1.pcpi_mul_rs1 [13]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_164 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_41 ), .B1
       (\genblk1.pcpi_mul_rs2 [19]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_759 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48949 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_198 ), .A1
       (\genblk1.pcpi_mul_rs1 [10]), .B0 (\genblk1.pcpi_mul_rs2 [25]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_69 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_758 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48950 (.A0
       (\genblk1.pcpi_mul_rs1 [3]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ), .B0
       (\genblk1.pcpi_mul_rs2 [11]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_93 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_757 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48951 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_197 ), .A1
       (\genblk1.pcpi_mul_rs1 [15]), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_97 ), .B1
       (\genblk1.pcpi_mul_rs2 [29]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_756 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48952 (.A0
       (\genblk1.pcpi_mul_rs1 [11]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_165 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_51 ), .B1
       (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_755 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48953 (.A0
       (\genblk1.pcpi_mul_rs1 [25]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_53 ), .B1
       (\genblk1.pcpi_mul_rs2 [11]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_754 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48954 (.A0
       (\genblk1.pcpi_mul_rs1 [24]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_166 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_99 ), .B1
       (\genblk1.pcpi_mul_rs2 [15]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_753 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48955 (.A0
       (\genblk1.pcpi_mul_rs1 [7]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_166 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_91 ), .B1
       (\genblk1.pcpi_mul_rs2 [15]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_752 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48956 (.A0
       (\genblk1.pcpi_mul_rs1 [18]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_79 ), .B1
       (\genblk1.pcpi_mul_rs2 [23]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_751 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48957 (.A0
       (\genblk1.pcpi_mul_rs1 [31]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_196 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_43 ), .B1
       (\genblk1.pcpi_mul_rs2 [13]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_750 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48958 (.A0
       (\genblk1.pcpi_mul_rs1 [29]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_195 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_61 ), .B1
       (\genblk1.pcpi_mul_rs2 [21]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_749 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48959 (.A0
       (\genblk1.pcpi_mul_rs1 [6]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_167 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_59 ), .B1
       (\genblk1.pcpi_mul_rs2 [7]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_748 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48960 (.A0
       (\genblk1.pcpi_mul_rs1 [8]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_170 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_85 ), .B1
       (\genblk1.pcpi_mul_rs2 [5]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_747 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48961 (.A0
       (\genblk1.pcpi_mul_rs1 [5]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_196 ), .B0
       (\genblk1.pcpi_mul_rs2 [13]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_47 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_746 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48962 (.A0
       (\genblk1.pcpi_mul_rs1 [16]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_195 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_89 ), .B1
       (\genblk1.pcpi_mul_rs2 [21]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_745 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48963 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ), .A1
       (\genblk1.pcpi_mul_rs1 [8]), .B0 (\genblk1.pcpi_mul_rs2 [23]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_85 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_744 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48964 (.A0
       (\genblk1.pcpi_mul_rs1 [18]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_195 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_79 ), .B1
       (\genblk1.pcpi_mul_rs2 [21]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_743 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48965 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_198 ), .A1
       (\genblk1.pcpi_mul_rs1 [16]), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_89 ), .B1
       (\genblk1.pcpi_mul_rs2 [25]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_742 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48966 (.A0
       (\genblk1.pcpi_mul_rs1 [26]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_193 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_55 ), .B1
       (\genblk1.pcpi_mul_rs2 [27]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_741 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48967 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_193 ), .A1
       (\genblk1.pcpi_mul_rs1 [5]), .B0 (\genblk1.pcpi_mul_rs2 [27]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_47 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_740 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48968 (.A0
       (\genblk1.pcpi_mul_rs1 [14]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_39 ), .B1
       (\genblk1.pcpi_mul_rs2 [11]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_739 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48969 (.A0
       (\genblk1.pcpi_mul_rs1 [18]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_196 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_79 ), .B1
       (\genblk1.pcpi_mul_rs2 [13]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_738 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48970 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_193 ), .A1
       (\genblk1.pcpi_mul_rs1 [9]), .B0 (\genblk1.pcpi_mul_rs2 [27]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_75 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_737 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48971 (.A0
       (\genblk1.pcpi_mul_rs1 [14]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_196 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_39 ), .B1
       (\genblk1.pcpi_mul_rs2 [13]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_736 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48972 (.A0
       (\genblk1.pcpi_mul_rs1 [16]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_166 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_89 ), .B1
       (\genblk1.pcpi_mul_rs2 [15]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_735 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48973 (.A0
       (\genblk1.pcpi_mul_rs1 [26]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_195 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_55 ), .B1
       (\genblk1.pcpi_mul_rs2 [21]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_734 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48974 (.A0
       (\genblk1.pcpi_mul_rs1 [17]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_193 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_83 ), .B1
       (\genblk1.pcpi_mul_rs2 [27]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_733 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48975 (.A0
       (\genblk1.pcpi_mul_rs1 [18]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_166 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_79 ), .B1
       (\genblk1.pcpi_mul_rs2 [15]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_732 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48976 (.A0
       (\genblk1.pcpi_mul_rs1 [1]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_170 ), .B0
       (\genblk1.pcpi_mul_rs2 [5]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_81 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_731 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48977 (.A0
       (\genblk1.pcpi_mul_rs1 [11]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_163 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_51 ), .B1
       (\genblk1.pcpi_mul_rs2 [9]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_730 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48978 (.A0
       (\genblk1.pcpi_mul_rs1 [16]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_194 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_89 ), .B1
       (\genblk1.pcpi_mul_rs2 [17]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_729 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48979 (.A0
       (\genblk1.pcpi_mul_rs1 [31]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_163 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_43 ), .B1
       (\genblk1.pcpi_mul_rs2 [9]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_728 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48980 (.A0
       (\genblk1.pcpi_mul_rs1 [28]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_165 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_65 ), .B1
       (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_727 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48981 (.A0
       (\genblk1.pcpi_mul_rs1 [27]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_196 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_77 ), .B1
       (\genblk1.pcpi_mul_rs2 [13]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_726 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48982 (.A0
       (\genblk1.pcpi_mul_rs1 [10]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_163 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_69 ), .B1
       (\genblk1.pcpi_mul_rs2 [9]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_725 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48983 (.A0
       (\genblk1.pcpi_mul_rs1 [22]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_163 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_95 ), .B1
       (\genblk1.pcpi_mul_rs2 [9]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_724 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48984 (.A0
       (\genblk1.pcpi_mul_rs1 [31]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_197 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_43 ), .B1
       (\genblk1.pcpi_mul_rs2 [29]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_723 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48985 (.A0
       (\genblk1.pcpi_mul_rs1 [22]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_164 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_95 ), .B1
       (\genblk1.pcpi_mul_rs2 [19]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_722 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48986 (.A0
       (\genblk1.pcpi_mul_rs1 [21]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_164 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_67 ), .B1
       (\genblk1.pcpi_mul_rs2 [19]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_721 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48987 (.A0
       (\genblk1.pcpi_mul_rs1 [29]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_198 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_61 ), .B1
       (\genblk1.pcpi_mul_rs2 [25]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_720 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48988 (.A0
       (\genblk1.pcpi_mul_rs1 [27]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_165 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_77 ), .B1
       (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_719 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48989 (.A0
       (\genblk1.pcpi_mul_rs1 [15]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_166 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_97 ), .B1
       (\genblk1.pcpi_mul_rs2 [15]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_718 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48990 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_198 ), .A1
       (\genblk1.pcpi_mul_rs1 [7]), .B0 (\genblk1.pcpi_mul_rs2 [25]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_91 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_717 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48991 (.A0
       (\genblk1.pcpi_mul_rs1 [16]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_165 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_89 ), .B1
       (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_716 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48992 (.A0
       (\genblk1.pcpi_mul_rs1 [29]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_61 ), .B1
       (\genblk1.pcpi_mul_rs2 [11]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_715 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48993 (.A0
       (\genblk1.pcpi_mul_rs1 [27]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_166 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_77 ), .B1
       (\genblk1.pcpi_mul_rs2 [15]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_714 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48994 (.A0
       (\genblk1.pcpi_mul_rs1 [24]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_163 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_99 ), .B1
       (\genblk1.pcpi_mul_rs2 [9]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_713 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48995 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ), .A1
       (\genblk1.pcpi_mul_rs1 [9]), .B0 (\genblk1.pcpi_mul_rs2 [23]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_75 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_712 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48996 (.A0
       (\genblk1.pcpi_mul_rs1 [19]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_163 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_73 ), .B1
       (\genblk1.pcpi_mul_rs2 [9]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_711 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48997 (.A0
       (\genblk1.pcpi_mul_rs1 [4]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ), .B0
       (\genblk1.pcpi_mul_rs2 [11]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_71 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_710 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48998 (.A0
       (\genblk1.pcpi_mul_rs1 [11]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_164 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_51 ), .B1
       (\genblk1.pcpi_mul_rs2 [19]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_709 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g48999 (.A0
       (\genblk1.pcpi_mul_rs1 [23]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_170 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_49 ), .B1
       (\genblk1.pcpi_mul_rs2 [5]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_708 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49000 (.A0
       (\genblk1.pcpi_mul_rs1 [22]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_197 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_95 ), .B1
       (\genblk1.pcpi_mul_rs2 [29]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_707 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49001 (.A0
       (\genblk1.pcpi_mul_rs1 [25]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_170 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_53 ), .B1
       (\genblk1.pcpi_mul_rs2 [5]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_706 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49002 (.A0
       (\genblk1.pcpi_mul_rs1 [19]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_197 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_73 ), .B1
       (\genblk1.pcpi_mul_rs2 [29]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_705 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49003 (.A0
       (\genblk1.pcpi_mul_rs1 [31]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_43 ), .B1
       (\genblk1.pcpi_mul_rs2 [23]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_704 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49004 (.A0
       (\genblk1.pcpi_mul_rs1 [19]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_73 ), .B1
       (\genblk1.pcpi_mul_rs2 [11]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_703 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49005 (.A0
       (\genblk1.pcpi_mul_rs1 [21]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_193 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_67 ), .B1
       (\genblk1.pcpi_mul_rs2 [27]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_702 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49006 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_197 ), .A1
       (\genblk1.pcpi_mul_rs1 [7]), .B0 (\genblk1.pcpi_mul_rs2 [29]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_91 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_701 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49007 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_198 ), .A1
       (\genblk1.pcpi_mul_rs1 [5]), .B0 (\genblk1.pcpi_mul_rs2 [25]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_47 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_700 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49008 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_193 ), .A1
       (\genblk1.pcpi_mul_rs1 [4]), .B0 (\genblk1.pcpi_mul_rs2 [27]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_71 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_699 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49009 (.A0
       (\genblk1.pcpi_mul_rs1 [29]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_193 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_61 ), .B1
       (\genblk1.pcpi_mul_rs2 [27]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_698 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49010 (.A0
       (\genblk1.pcpi_mul_rs1 [25]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_197 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_53 ), .B1
       (\genblk1.pcpi_mul_rs2 [29]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_697 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49011 (.A0
       (\genblk1.pcpi_mul_rs1 [25]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_164 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_53 ), .B1
       (\genblk1.pcpi_mul_rs2 [19]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_696 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49012 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_164 ), .A1
       (\genblk1.pcpi_mul_rs1 [4]), .B0 (\genblk1.pcpi_mul_rs2 [19]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_71 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_695 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49013 (.A0
       (\genblk1.pcpi_mul_rs1 [28]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_193 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_65 ), .B1
       (\genblk1.pcpi_mul_rs2 [27]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_694 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49014 (.A0
       (\genblk1.pcpi_mul_rs1 [23]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_165 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_49 ), .B1
       (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_693 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49015 (.A0
       (\genblk1.pcpi_mul_rs1 [28]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_198 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_65 ), .B1
       (\genblk1.pcpi_mul_rs2 [25]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_692 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49016 (.A0
       (\genblk1.pcpi_mul_rs1 [12]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_196 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_45 ), .B1
       (\genblk1.pcpi_mul_rs2 [13]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_691 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49017 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_195 ), .A1
       (\genblk1.pcpi_mul_rs1 [8]), .B0 (\genblk1.pcpi_mul_rs2 [21]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_85 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_690 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49018 (.A0
       (\genblk1.pcpi_mul_rs1 [18]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_163 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_79 ), .B1
       (\genblk1.pcpi_mul_rs2 [9]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_689 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49019 (.A0
       (\genblk1.pcpi_mul_rs1 [24]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_170 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_99 ), .B1
       (\genblk1.pcpi_mul_rs2 [5]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_688 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49020 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_193 ), .A1
       (\genblk1.pcpi_mul_rs1 [11]), .B0 (\genblk1.pcpi_mul_rs2 [27]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_51 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_687 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49021 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_198 ), .A1
       (\genblk1.pcpi_mul_rs1 [4]), .B0 (\genblk1.pcpi_mul_rs2 [25]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_71 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_686 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49022 (.A0
       (\genblk1.pcpi_mul_rs1 [16]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_196 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_89 ), .B1
       (\genblk1.pcpi_mul_rs2 [13]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_685 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49023 (.A0
       (\genblk1.pcpi_mul_rs1 [31]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_198 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_43 ), .B1
       (\genblk1.pcpi_mul_rs2 [25]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_684 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49024 (.A0
       (\genblk1.pcpi_mul_rs1 [16]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_89 ), .B1
       (\genblk1.pcpi_mul_rs2 [23]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_683 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49025 (.A0
       (\genblk1.pcpi_mul_rs1 [23]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_195 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_49 ), .B1
       (\genblk1.pcpi_mul_rs2 [21]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_682 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49026 (.A0
       (\genblk1.pcpi_mul_rs1 [20]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_196 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_87 ), .B1
       (\genblk1.pcpi_mul_rs2 [13]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_681 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49027 (.A0
       (\genblk1.pcpi_mul_rs1 [5]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_163 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_47 ), .B1
       (\genblk1.pcpi_mul_rs2 [9]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_680 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49028 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_197 ), .A1
       (\genblk1.pcpi_mul_rs1 [1]), .B0 (\genblk1.pcpi_mul_rs2 [29]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_81 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_679 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49029 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_193 ), .A1
       (\genblk1.pcpi_mul_rs1 [12]), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_45 ), .B1
       (\genblk1.pcpi_mul_rs2 [27]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_678 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49030 (.A0
       (\genblk1.pcpi_mul_rs1 [23]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_49 ), .B1
       (\genblk1.pcpi_mul_rs2 [23]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_677 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49031 (.A0
       (\genblk1.pcpi_mul_rs1 [26]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_165 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_55 ), .B1
       (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_676 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49032 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_193 ), .A1
       (\genblk1.pcpi_mul_rs1 [13]), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_41 ), .B1
       (\genblk1.pcpi_mul_rs2 [27]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_675 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49033 (.A0
       (\genblk1.pcpi_mul_rs1 [6]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_59 ), .B1
       (\genblk1.pcpi_mul_rs2 [11]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_674 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49034 (.A0
       (\genblk1.pcpi_mul_rs1 [26]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_196 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_55 ), .B1
       (\genblk1.pcpi_mul_rs2 [13]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_673 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49035 (.A0
       (\genblk1.pcpi_mul_rs1 [24]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_195 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_99 ), .B1
       (\genblk1.pcpi_mul_rs2 [21]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_672 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49036 (.A0
       (\genblk1.pcpi_mul_rs1 [14]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_166 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_39 ), .B1
       (\genblk1.pcpi_mul_rs2 [15]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_671 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49037 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_195 ), .A1
       (\genblk1.pcpi_mul_rs1 [4]), .B0 (\genblk1.pcpi_mul_rs2 [21]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_71 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_670 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49038 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_193 ), .A1
       (\genblk1.pcpi_mul_rs1 [2]), .B0 (\genblk1.pcpi_mul_rs2 [27]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_57 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_669 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49039 (.A0
       (\genblk1.pcpi_mul_rs1 [4]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_170 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_71 ), .B1
       (\genblk1.pcpi_mul_rs2 [5]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_668 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49040 (.A0
       (\genblk1.pcpi_mul_rs1 [23]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_194 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_49 ), .B1
       (\genblk1.pcpi_mul_rs2 [17]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_667 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49041 (.A0
       (\genblk1.pcpi_mul_rs1 [28]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_166 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_65 ), .B1
       (\genblk1.pcpi_mul_rs2 [15]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_666 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49042 (.A0
       (\genblk1.pcpi_mul_rs1 [6]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_165 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_59 ), .B1
       (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_665 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49043 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_195 ), .A1
       (\genblk1.pcpi_mul_rs1 [17]), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_83 ), .B1
       (\genblk1.pcpi_mul_rs2 [21]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_664 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49044 (.A0
       (\genblk1.pcpi_mul_rs1 [16]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_89 ), .B1
       (\genblk1.pcpi_mul_rs2 [11]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_663 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49045 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_195 ), .A1
       (\genblk1.pcpi_mul_rs1 [14]), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_39 ), .B1
       (\genblk1.pcpi_mul_rs2 [21]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_662 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49046 (.A0
       (\genblk1.pcpi_mul_rs1 [28]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_164 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_65 ), .B1
       (\genblk1.pcpi_mul_rs2 [19]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_661 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49047 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_197 ), .A1
       (\genblk1.pcpi_mul_rs1 [18]), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_79 ), .B1
       (\genblk1.pcpi_mul_rs2 [29]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_660 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49048 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_193 ), .A1
       (\genblk1.pcpi_mul_rs1 [16]), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_89 ), .B1
       (\genblk1.pcpi_mul_rs2 [27]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_659 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49049 (.A0
       (\genblk1.pcpi_mul_rs1 [28]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_170 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_65 ), .B1
       (\genblk1.pcpi_mul_rs2 [5]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_658 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49050 (.A0
       (\genblk1.pcpi_mul_rs1 [25]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_198 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_53 ), .B1
       (\genblk1.pcpi_mul_rs2 [25]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_657 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49051 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_193 ), .A1
       (\genblk1.pcpi_mul_rs1 [6]), .B0 (\genblk1.pcpi_mul_rs2 [27]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_59 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_656 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49052 (.A0
       (\genblk1.pcpi_mul_rs1 [11]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_194 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_51 ), .B1
       (\genblk1.pcpi_mul_rs2 [17]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_655 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49053 (.A0
       (\genblk1.pcpi_mul_rs1 [11]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_170 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_51 ), .B1
       (\genblk1.pcpi_mul_rs2 [5]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_654 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49054 (.A0
       (\genblk1.pcpi_mul_rs1 [13]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_170 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_41 ), .B1
       (\genblk1.pcpi_mul_rs2 [5]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_653 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49055 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_193 ), .A1
       (\genblk1.pcpi_mul_rs1 [15]), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_97 ), .B1
       (\genblk1.pcpi_mul_rs2 [27]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_652 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49056 (.A0
       (\genblk1.pcpi_mul_rs1 [12]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_165 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_45 ), .B1
       (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_651 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49057 (.A0
       (\genblk1.pcpi_mul_rs1 [24]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_167 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_99 ), .B1
       (\genblk1.pcpi_mul_rs2 [7]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_650 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49058 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_193 ), .A1
       (\genblk1.pcpi_mul_rs1 [10]), .B0 (\genblk1.pcpi_mul_rs2 [27]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_69 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_649 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49059 (.A0
       (\genblk1.pcpi_mul_rs1 [23]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_197 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_49 ), .B1
       (\genblk1.pcpi_mul_rs2 [29]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_648 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49060 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ), .A1
       (\genblk1.pcpi_mul_rs1 [7]), .B0 (\genblk1.pcpi_mul_rs2 [23]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_91 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_647 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49061 (.A0
       (\genblk1.pcpi_mul_rs1 [9]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_164 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_75 ), .B1
       (\genblk1.pcpi_mul_rs2 [19]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_646 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49062 (.A0
       (\genblk1.pcpi_mul_rs1 [15]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_97 ), .B1
       (\genblk1.pcpi_mul_rs2 [23]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_645 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49063 (.A0
       (\genblk1.pcpi_mul_rs1 [5]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_170 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_47 ), .B1
       (\genblk1.pcpi_mul_rs2 [5]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_644 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49064 (.A0
       (\genblk1.pcpi_mul_rs1 [2]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_165 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_57 ), .B1
       (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_643 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49065 (.A0
       (\genblk1.pcpi_mul_rs1 [11]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_51 ), .B1
       (\genblk1.pcpi_mul_rs2 [11]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_642 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49066 (.A0
       (\genblk1.pcpi_mul_rs1 [25]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_196 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_53 ), .B1
       (\genblk1.pcpi_mul_rs2 [13]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_641 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49067 (.A0
       (\genblk1.pcpi_mul_rs1 [10]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_69 ), .B1
       (\genblk1.pcpi_mul_rs2 [11]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_640 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49068 (.A0
       (\genblk1.pcpi_mul_rs1 [20]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_195 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_87 ), .B1
       (\genblk1.pcpi_mul_rs2 [21]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_639 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49069 (.A0
       (\genblk1.pcpi_mul_rs1 [3]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_170 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_93 ), .B1
       (\genblk1.pcpi_mul_rs2 [5]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_638 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49070 (.A0
       (\genblk1.pcpi_mul_rs1 [27]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_77 ), .B1
       (\genblk1.pcpi_mul_rs2 [11]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_637 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49071 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_198 ), .A1
       (\genblk1.pcpi_mul_rs1 [3]), .B0 (\genblk1.pcpi_mul_rs2 [25]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_93 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_636 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49072 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_197 ), .A1
       (\genblk1.pcpi_mul_rs1 [9]), .B0 (\genblk1.pcpi_mul_rs2 [29]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_75 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_635 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49073 (.A0
       (\genblk1.pcpi_mul_rs1 [15]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_196 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_97 ), .B1
       (\genblk1.pcpi_mul_rs2 [13]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_634 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49074 (.A0
       (\genblk1.pcpi_mul_rs1 [21]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_166 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_67 ), .B1
       (\genblk1.pcpi_mul_rs2 [15]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_633 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49075 (.A0
       (\genblk1.pcpi_mul_rs1 [23]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_193 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_49 ), .B1
       (\genblk1.pcpi_mul_rs2 [27]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_632 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49076 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ), .A1
       (\genblk1.pcpi_mul_rs1 [4]), .B0 (\genblk1.pcpi_mul_rs2 [23]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_71 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_631 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49077 (.A0
       (\genblk1.pcpi_mul_rs1 [23]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_166 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_49 ), .B1
       (\genblk1.pcpi_mul_rs2 [15]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_630 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49078 (.A0
       (\genblk1.pcpi_mul_rs1 [27]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_195 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_77 ), .B1
       (\genblk1.pcpi_mul_rs2 [21]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_629 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49079 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_198 ), .A1
       (\genblk1.pcpi_mul_rs1 [14]), .B0 (\genblk1.pcpi_mul_rs2 [25]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_39 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_628 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49080 (.A0
       (\genblk1.pcpi_mul_rs1 [20]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_193 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_87 ), .B1
       (\genblk1.pcpi_mul_rs2 [27]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_627 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49081 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ), .A1
       (\genblk1.pcpi_mul_rs1 [6]), .B0 (\genblk1.pcpi_mul_rs2 [23]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_59 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_626 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49082 (.A0
       (\genblk1.pcpi_mul_rs1 [15]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_165 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_97 ), .B1
       (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_625 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49083 (.A0
       (\genblk1.pcpi_mul_rs1 [22]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_198 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_95 ), .B1
       (\genblk1.pcpi_mul_rs2 [25]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_624 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49084 (.A0
       (\genblk1.pcpi_mul_rs1 [24]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_164 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_99 ), .B1
       (\genblk1.pcpi_mul_rs2 [19]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_623 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49085 (.A0
       (\genblk1.pcpi_mul_rs1 [27]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_197 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_77 ), .B1
       (\genblk1.pcpi_mul_rs2 [29]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_622 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49086 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_195 ), .A1
       (\genblk1.pcpi_mul_rs1 [6]), .B0 (\genblk1.pcpi_mul_rs2 [21]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_59 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_621 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49087 (.A0
       (\genblk1.pcpi_mul_rs1 [22]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_95 ), .B1
       (\genblk1.pcpi_mul_rs2 [11]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_620 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49088 (.A0
       (\genblk1.pcpi_mul_rs1 [10]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_167 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_69 ), .B1
       (\genblk1.pcpi_mul_rs2 [7]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_619 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49089 (.A0
       (\genblk1.pcpi_mul_rs1 [10]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_194 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_69 ), .B1
       (\genblk1.pcpi_mul_rs2 [17]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_618 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49090 (.A0
       (\genblk1.pcpi_mul_rs1 [25]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_195 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_53 ), .B1
       (\genblk1.pcpi_mul_rs2 [21]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_617 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49091 (.A0
       (\genblk1.pcpi_mul_rs1 [24]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_194 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_99 ), .B1
       (\genblk1.pcpi_mul_rs2 [17]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_616 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49092 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_193 ), .A1
       (\genblk1.pcpi_mul_rs1 [8]), .B0 (\genblk1.pcpi_mul_rs2 [27]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_85 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_615 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49093 (.A0
       (\genblk1.pcpi_mul_rs1 [13]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_196 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_41 ), .B1
       (\genblk1.pcpi_mul_rs2 [13]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_614 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49094 (.A0
       (\genblk1.pcpi_mul_rs1 [29]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_165 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_61 ), .B1
       (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_613 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49095 (.A0
       (\genblk1.pcpi_mul_rs1 [9]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_75 ), .B1
       (\genblk1.pcpi_mul_rs2 [11]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_612 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49096 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_194 ), .A1
       (\genblk1.pcpi_mul_rs1 [1]), .B0 (\genblk1.pcpi_mul_rs2 [17]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_81 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_611 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49097 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_193 ), .A1
       (\genblk1.pcpi_mul_rs1 [7]), .B0 (\genblk1.pcpi_mul_rs2 [27]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_91 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_610 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49098 (.A0
       (\genblk1.pcpi_mul_rs1 [2]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_167 ), .B0
       (\genblk1.pcpi_mul_rs2 [7]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_57 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_609 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49099 (.A0
       (\genblk1.pcpi_mul_rs1 [19]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_195 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_73 ), .B1
       (\genblk1.pcpi_mul_rs2 [21]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_608 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49100 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_193 ), .A1
       (\genblk1.pcpi_mul_rs1 [14]), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_39 ), .B1
       (\genblk1.pcpi_mul_rs2 [27]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_607 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49101 (.A0
       (\genblk1.pcpi_mul_rs1 [27]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_167 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_77 ), .B1
       (\genblk1.pcpi_mul_rs2 [7]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_606 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49102 (.A0
       (\genblk1.pcpi_mul_rs1 [13]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_165 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_41 ), .B1
       (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_605 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49103 (.A0
       (\genblk1.pcpi_mul_rs1 [13]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_195 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_41 ), .B1
       (\genblk1.pcpi_mul_rs2 [21]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_604 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49104 (.A0
       (\genblk1.pcpi_mul_rs1 [21]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_196 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_67 ), .B1
       (\genblk1.pcpi_mul_rs2 [13]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_603 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49105 (.A0
       (\genblk1.pcpi_mul_rs1 [30]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_197 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_63 ), .B1
       (\genblk1.pcpi_mul_rs2 [29]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_602 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49106 (.A0
       (\genblk1.pcpi_mul_rs1 [9]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_170 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_75 ), .B1
       (\genblk1.pcpi_mul_rs2 [5]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_601 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49107 (.A0
       (\genblk1.pcpi_mul_rs1 [18]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_79 ), .B1
       (\genblk1.pcpi_mul_rs2 [11]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_600 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49108 (.A0
       (\genblk1.pcpi_mul_rs1 [20]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_167 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_87 ), .B1
       (\genblk1.pcpi_mul_rs2 [7]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_599 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49109 (.A0
       (\genblk1.pcpi_mul_rs1 [7]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_194 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_91 ), .B1
       (\genblk1.pcpi_mul_rs2 [17]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_598 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49110 (.A0
       (\genblk1.pcpi_mul_rs1 [19]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_167 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_73 ), .B1
       (\genblk1.pcpi_mul_rs2 [7]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_597 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49111 (.A0
       (\genblk1.pcpi_mul_rs1 [24]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_197 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_99 ), .B1
       (\genblk1.pcpi_mul_rs2 [29]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_596 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49112 (.A0
       (\genblk1.pcpi_mul_rs1 [19]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_193 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_73 ), .B1
       (\genblk1.pcpi_mul_rs2 [27]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_595 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49113 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_194 ), .A1
       (\genblk1.pcpi_mul_rs1 [3]), .B0 (\genblk1.pcpi_mul_rs2 [17]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_93 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_594 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49114 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_195 ), .A1
       (\genblk1.pcpi_mul_rs1 [5]), .B0 (\genblk1.pcpi_mul_rs2 [21]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_47 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_593 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49115 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_197 ), .A1
       (\genblk1.pcpi_mul_rs1 [12]), .B0 (\genblk1.pcpi_mul_rs2 [29]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_45 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_592 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49116 (.A0
       (\genblk1.pcpi_mul_rs1 [5]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_164 ), .B0
       (\genblk1.pcpi_mul_rs2 [19]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_47 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_591 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49117 (.A0
       (\genblk1.pcpi_mul_rs1 [10]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_196 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_69 ), .B1
       (\genblk1.pcpi_mul_rs2 [13]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_590 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49118 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_198 ), .A1
       (\genblk1.pcpi_mul_rs1 [1]), .B0 (\genblk1.pcpi_mul_rs2 [25]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_81 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_589 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49119 (.A0
       (\genblk1.pcpi_mul_rs1 [12]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_163 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_45 ), .B1
       (\genblk1.pcpi_mul_rs2 [9]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_588 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49120 (.A0
       (\genblk1.pcpi_mul_rs1 [11]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_166 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_51 ), .B1
       (\genblk1.pcpi_mul_rs2 [15]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_587 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49121 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_195 ), .A1
       (\genblk1.pcpi_mul_rs1 [9]), .B0 (\genblk1.pcpi_mul_rs2 [21]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_75 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_586 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49122 (.A0
       (\genblk1.pcpi_mul_rs1 [23]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_198 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_49 ), .B1
       (\genblk1.pcpi_mul_rs2 [25]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_585 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49123 (.A0
       (\genblk1.pcpi_mul_rs1 [12]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_166 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_45 ), .B1
       (\genblk1.pcpi_mul_rs2 [15]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_584 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49124 (.A0
       (\genblk1.pcpi_mul_rs1 [22]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_193 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_95 ), .B1
       (\genblk1.pcpi_mul_rs2 [27]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_583 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49125 (.A0
       (\genblk1.pcpi_mul_rs1 [22]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_195 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_95 ), .B1
       (\genblk1.pcpi_mul_rs2 [21]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_582 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49126 (.A0
       (\genblk1.pcpi_mul_rs1 [15]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_97 ), .B1
       (\genblk1.pcpi_mul_rs2 [11]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_581 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49127 (.A0
       (\genblk1.pcpi_mul_rs1 [19]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_196 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_73 ), .B1
       (\genblk1.pcpi_mul_rs2 [13]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_580 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49128 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_194 ), .A1
       (\genblk1.pcpi_mul_rs1 [4]), .B0 (\genblk1.pcpi_mul_rs2 [17]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_71 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_579 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49129 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_195 ), .A1
       (\genblk1.pcpi_mul_rs1 [10]), .B0 (\genblk1.pcpi_mul_rs2 [21]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_69 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_578 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49130 (.A0
       (\genblk1.pcpi_mul_rs1 [24]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_165 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_99 ), .B1
       (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_577 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49131 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_195 ), .A1
       (\genblk1.pcpi_mul_rs1 [1]), .B0 (\genblk1.pcpi_mul_rs2 [21]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_81 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_576 ));
  AND2X2 \genblk1.pcpi_mul_mul_2366_47_g49132 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_221 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_226 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_137 ));
  XNOR2X2 \genblk1.pcpi_mul_mul_2366_47_g49133 (.A
       (\genblk1.pcpi_mul_rs2 [26]), .B (\genblk1.pcpi_mul_rs2 [25]),
       .Y (\genblk1.pcpi_mul_mul_2366_47_n_574 ));
  XNOR2X2 \genblk1.pcpi_mul_mul_2366_47_g49134 (.A
       (\genblk1.pcpi_mul_rs2 [10]), .B (\genblk1.pcpi_mul_rs2 [9]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ));
  XNOR2X2 \genblk1.pcpi_mul_mul_2366_47_g49135 (.A
       (\genblk1.pcpi_mul_rs2 [4]), .B (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ));
  XNOR2X2 \genblk1.pcpi_mul_mul_2366_47_g49136 (.A
       (\genblk1.pcpi_mul_rs2 [16]), .B (\genblk1.pcpi_mul_rs2 [15]),
       .Y (\genblk1.pcpi_mul_mul_2366_47_n_571 ));
  XNOR2X2 \genblk1.pcpi_mul_mul_2366_47_g49137 (.A
       (\genblk1.pcpi_mul_rs2 [24]), .B (\genblk1.pcpi_mul_rs2 [23]),
       .Y (\genblk1.pcpi_mul_mul_2366_47_n_570 ));
  XNOR2X2 \genblk1.pcpi_mul_mul_2366_47_g49138 (.A
       (\genblk1.pcpi_mul_rs2 [30]), .B (\genblk1.pcpi_mul_rs2 [29]),
       .Y (\genblk1.pcpi_mul_mul_2366_47_n_569 ));
  XNOR2X2 \genblk1.pcpi_mul_mul_2366_47_g49139 (.A
       (\genblk1.pcpi_mul_rs2 [6]), .B (\genblk1.pcpi_mul_rs2 [5]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ));
  XNOR2X2 \genblk1.pcpi_mul_mul_2366_47_g49140 (.A
       (\genblk1.pcpi_mul_rs2 [18]), .B (\genblk1.pcpi_mul_rs2 [17]),
       .Y (\genblk1.pcpi_mul_mul_2366_47_n_567 ));
  XNOR2X2 \genblk1.pcpi_mul_mul_2366_47_g49141 (.A
       (\genblk1.pcpi_mul_rs2 [8]), .B (\genblk1.pcpi_mul_rs2 [7]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ));
  XNOR2X2 \genblk1.pcpi_mul_mul_2366_47_g49142 (.A
       (\genblk1.pcpi_mul_rs2 [20]), .B (\genblk1.pcpi_mul_rs2 [19]),
       .Y (\genblk1.pcpi_mul_mul_2366_47_n_565 ));
  XNOR2X2 \genblk1.pcpi_mul_mul_2366_47_g49143 (.A
       (\genblk1.pcpi_mul_rs2 [14]), .B (\genblk1.pcpi_mul_rs2 [13]),
       .Y (\genblk1.pcpi_mul_mul_2366_47_n_564 ));
  XNOR2X2 \genblk1.pcpi_mul_mul_2366_47_g49144 (.A
       (\genblk1.pcpi_mul_rs2 [22]), .B (\genblk1.pcpi_mul_rs2 [21]),
       .Y (\genblk1.pcpi_mul_mul_2366_47_n_563 ));
  XNOR2X2 \genblk1.pcpi_mul_mul_2366_47_g49145 (.A
       (\genblk1.pcpi_mul_rs2 [28]), .B (\genblk1.pcpi_mul_rs2 [27]),
       .Y (\genblk1.pcpi_mul_mul_2366_47_n_562 ));
  XNOR2X2 \genblk1.pcpi_mul_mul_2366_47_g49146 (.A
       (\genblk1.pcpi_mul_rs2 [2]), .B (\genblk1.pcpi_mul_rs2 [1]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ));
  XNOR2X2 \genblk1.pcpi_mul_mul_2366_47_g49147 (.A
       (\genblk1.pcpi_mul_rs2 [12]), .B (\genblk1.pcpi_mul_rs2 [11]),
       .Y (\genblk1.pcpi_mul_mul_2366_47_n_560 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_g49148 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_345 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_346 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_g49149 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_341 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_342 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_g49150 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_338 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_339 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_g49151 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_334 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_335 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_g49152 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_327 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_328 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_g49153 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_324 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_325 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_g49154 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_320 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_321 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_g49155 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_318 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_319 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_g49156 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_313 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_314 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_g49157 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_305 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_306 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_g49158 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_298 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_299 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_g49159 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_293 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_294 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_g49160 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_289 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_290 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_g49161 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_286 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_287 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_g49162 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_281 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_282 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_g49163 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_279 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_280 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_g49164 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_276 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_277 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_g49165 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_273 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_274 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_g49166 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_270 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_271 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49167 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ), .A1
       (\genblk1.pcpi_mul_rs1 [0]), .B0 (\genblk1.pcpi_mul_rs2 [11]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_251 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g49168 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .A1
       (\genblk1.pcpi_mul_rs2 [1]), .B0 (\genblk1.pcpi_mul_rs1 [0]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_171 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_250 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49169 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_167 ), .A1
       (\genblk1.pcpi_mul_rs1 [0]), .B0 (\genblk1.pcpi_mul_rs2 [7]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_249 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49170 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_198 ), .A1
       (\genblk1.pcpi_mul_rs1 [0]), .B0 (\genblk1.pcpi_mul_rs2 [25]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_248 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49171 (.A0
       (\genblk1.pcpi_mul_rs1 [0]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_165 ), .B0
       (\genblk1.pcpi_mul_rs2 [3]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_247 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49172 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_164 ), .A1
       (\genblk1.pcpi_mul_rs1 [0]), .B0 (\genblk1.pcpi_mul_rs2 [19]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_246 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49173 (.A0
       (\genblk1.pcpi_mul_rs1 [0]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_170 ), .B0
       (\genblk1.pcpi_mul_rs2 [5]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_245 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49174 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_197 ), .A1
       (\genblk1.pcpi_mul_rs1 [0]), .B0 (\genblk1.pcpi_mul_rs2 [29]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_244 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49175 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_163 ), .A1
       (\genblk1.pcpi_mul_rs1 [0]), .B0 (\genblk1.pcpi_mul_rs2 [9]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_243 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49176 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_195 ), .A1
       (\genblk1.pcpi_mul_rs1 [0]), .B0 (\genblk1.pcpi_mul_rs2 [21]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_242 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49177 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_196 ), .A1
       (\genblk1.pcpi_mul_rs1 [0]), .B0 (\genblk1.pcpi_mul_rs2 [13]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_241 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49178 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_166 ), .A1
       (\genblk1.pcpi_mul_rs1 [0]), .B0 (\genblk1.pcpi_mul_rs2 [15]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_240 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49179 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ), .A1
       (\genblk1.pcpi_mul_rs1 [0]), .B0 (\genblk1.pcpi_mul_rs2 [23]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_239 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49180 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_194 ), .A1
       (\genblk1.pcpi_mul_rs1 [0]), .B0 (\genblk1.pcpi_mul_rs2 [17]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_238 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49181 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_193 ), .A1
       (\genblk1.pcpi_mul_rs1 [0]), .B0 (\genblk1.pcpi_mul_rs2 [27]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_237 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49182 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .A1
       (\genblk1.pcpi_mul_rs1 [0]), .B0 (\genblk1.pcpi_mul_rs2 [31]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_236 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49183 (.A0
       (\genblk1.pcpi_mul_rs1 [30]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_63 ), .B1
       (\genblk1.pcpi_mul_rs2 [23]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_537 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49184 (.A0
       (\genblk1.pcpi_mul_rs1 [18]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_193 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_79 ), .B1
       (\genblk1.pcpi_mul_rs2 [27]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_536 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49185 (.A0
       (\genblk1.pcpi_mul_rs1 [31]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_193 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_43 ), .B1
       (\genblk1.pcpi_mul_rs2 [27]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_535 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49186 (.A0
       (\genblk1.pcpi_mul_rs1 [25]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_165 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_53 ), .B1
       (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_534 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49187 (.A0
       (\genblk1.pcpi_mul_rs1 [30]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_170 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_63 ), .B1
       (\genblk1.pcpi_mul_rs2 [5]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_533 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49188 (.A0
       (\genblk1.pcpi_mul_rs1 [21]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_163 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_67 ), .B1
       (\genblk1.pcpi_mul_rs2 [9]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_532 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49189 (.A0
       (\genblk1.pcpi_mul_rs1 [21]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_167 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_67 ), .B1
       (\genblk1.pcpi_mul_rs2 [7]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_531 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49190 (.A0
       (\genblk1.pcpi_mul_rs1 [16]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_163 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_89 ), .B1
       (\genblk1.pcpi_mul_rs2 [9]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_530 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49191 (.A0
       (\genblk1.pcpi_mul_rs1 [19]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_165 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_73 ), .B1
       (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_529 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49192 (.A0
       (\genblk1.pcpi_mul_rs1 [26]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_55 ), .B1
       (\genblk1.pcpi_mul_rs2 [23]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_528 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49193 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_197 ), .A1
       (\genblk1.pcpi_mul_rs1 [5]), .B0 (\genblk1.pcpi_mul_rs2 [29]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_47 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_527 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49194 (.A0
       (\genblk1.pcpi_mul_rs1 [12]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_45 ), .B1
       (\genblk1.pcpi_mul_rs2 [11]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_526 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49195 (.A0
       (\genblk1.pcpi_mul_rs1 [15]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_164 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_97 ), .B1
       (\genblk1.pcpi_mul_rs2 [19]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_525 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49196 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_197 ), .A1
       (\genblk1.pcpi_mul_rs1 [4]), .B0 (\genblk1.pcpi_mul_rs2 [29]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_71 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_524 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49197 (.A0
       (\genblk1.pcpi_mul_rs1 [9]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_196 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_75 ), .B1
       (\genblk1.pcpi_mul_rs2 [13]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_523 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49198 (.A0
       (\genblk1.pcpi_mul_rs1 [6]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_170 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_59 ), .B1
       (\genblk1.pcpi_mul_rs2 [5]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_522 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49199 (.A0
       (\genblk1.pcpi_mul_rs1 [23]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_167 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_49 ), .B1
       (\genblk1.pcpi_mul_rs2 [7]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_521 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49200 (.A0
       (\genblk1.pcpi_mul_rs1 [8]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_166 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_85 ), .B1
       (\genblk1.pcpi_mul_rs2 [15]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_520 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49201 (.A0
       (\genblk1.pcpi_mul_rs1 [23]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_196 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_49 ), .B1
       (\genblk1.pcpi_mul_rs2 [13]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_519 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49202 (.A0
       (\genblk1.pcpi_mul_rs1 [17]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_165 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_83 ), .B1
       (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_518 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49203 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_196 ), .A1
       (\genblk1.pcpi_mul_rs1 [1]), .B0 (\genblk1.pcpi_mul_rs2 [13]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_81 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_517 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49204 (.A0
       (\genblk1.pcpi_mul_rs1 [26]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_164 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_55 ), .B1
       (\genblk1.pcpi_mul_rs2 [19]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_516 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49205 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_198 ), .A1
       (\genblk1.pcpi_mul_rs1 [6]), .B0 (\genblk1.pcpi_mul_rs2 [25]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_59 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_515 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49206 (.A0
       (\genblk1.pcpi_mul_rs1 [28]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_194 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_65 ), .B1
       (\genblk1.pcpi_mul_rs2 [17]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_514 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49207 (.A0
       (\genblk1.pcpi_mul_rs1 [20]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_197 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_87 ), .B1
       (\genblk1.pcpi_mul_rs2 [29]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_513 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49208 (.A0
       (\genblk1.pcpi_mul_rs1 [17]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_167 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_83 ), .B1
       (\genblk1.pcpi_mul_rs2 [7]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_512 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49209 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_195 ), .A1
       (\genblk1.pcpi_mul_rs1 [2]), .B0 (\genblk1.pcpi_mul_rs2 [21]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_57 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_511 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49210 (.A0
       (\genblk1.pcpi_mul_rs1 [3]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_166 ), .B0
       (\genblk1.pcpi_mul_rs2 [15]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_93 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_510 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49211 (.A0
       (\genblk1.pcpi_mul_rs1 [18]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_194 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_79 ), .B1
       (\genblk1.pcpi_mul_rs2 [17]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_509 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49212 (.A0
       (\genblk1.pcpi_mul_rs1 [26]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_198 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_55 ), .B1
       (\genblk1.pcpi_mul_rs2 [25]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_508 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49213 (.A0
       (\genblk1.pcpi_mul_rs1 [27]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_164 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_77 ), .B1
       (\genblk1.pcpi_mul_rs2 [19]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_507 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49214 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_164 ), .A1
       (\genblk1.pcpi_mul_rs1 [1]), .B0 (\genblk1.pcpi_mul_rs2 [19]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_81 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_506 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49215 (.A0
       (\genblk1.pcpi_mul_rs1 [2]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_163 ), .B0
       (\genblk1.pcpi_mul_rs2 [9]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_57 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_505 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49216 (.A0
       (\genblk1.pcpi_mul_rs1 [5]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_194 ), .B0
       (\genblk1.pcpi_mul_rs2 [17]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_47 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_504 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49217 (.A0
       (\genblk1.pcpi_mul_rs1 [21]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_165 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_67 ), .B1
       (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_503 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49218 (.A0
       (\genblk1.pcpi_mul_rs1 [21]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_194 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_67 ), .B1
       (\genblk1.pcpi_mul_rs2 [17]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_502 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49219 (.A0
       (\genblk1.pcpi_mul_rs1 [17]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_166 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_83 ), .B1
       (\genblk1.pcpi_mul_rs2 [15]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_501 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49220 (.A0
       (\genblk1.pcpi_mul_rs1 [30]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_166 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_63 ), .B1
       (\genblk1.pcpi_mul_rs2 [15]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_500 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49221 (.A0
       (\genblk1.pcpi_mul_rs1 [17]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_164 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_83 ), .B1
       (\genblk1.pcpi_mul_rs2 [19]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_499 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49222 (.A0
       (\genblk1.pcpi_mul_rs1 [16]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_164 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_89 ), .B1
       (\genblk1.pcpi_mul_rs2 [19]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_498 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49223 (.A0
       (\genblk1.pcpi_mul_rs1 [20]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_198 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_87 ), .B1
       (\genblk1.pcpi_mul_rs2 [25]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_497 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49224 (.A0
       (\genblk1.pcpi_mul_rs1 [30]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_198 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_63 ), .B1
       (\genblk1.pcpi_mul_rs2 [25]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_496 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49225 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_197 ), .A1
       (\genblk1.pcpi_mul_rs1 [10]), .B0 (\genblk1.pcpi_mul_rs2 [29]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_69 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_495 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49226 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_198 ), .A1
       (\genblk1.pcpi_mul_rs1 [19]), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_73 ), .B1
       (\genblk1.pcpi_mul_rs2 [25]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_494 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49227 (.A0
       (\genblk1.pcpi_mul_rs1 [13]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_163 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_41 ), .B1
       (\genblk1.pcpi_mul_rs2 [9]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_493 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49228 (.A0
       (\genblk1.pcpi_mul_rs1 [12]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_195 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_45 ), .B1
       (\genblk1.pcpi_mul_rs2 [21]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_492 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49229 (.A0
       (\genblk1.pcpi_mul_rs1 [29]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_166 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_61 ), .B1
       (\genblk1.pcpi_mul_rs2 [15]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_491 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49230 (.A0
       (\genblk1.pcpi_mul_rs1 [26]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_170 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_55 ), .B1
       (\genblk1.pcpi_mul_rs2 [5]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_490 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49231 (.A0
       (\genblk1.pcpi_mul_rs1 [24]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_99 ), .B1
       (\genblk1.pcpi_mul_rs2 [23]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_489 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49232 (.A0
       (\genblk1.pcpi_mul_rs1 [9]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_194 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_75 ), .B1
       (\genblk1.pcpi_mul_rs2 [17]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_488 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49233 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ), .A1
       (\genblk1.pcpi_mul_rs1 [10]), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_69 ), .B1
       (\genblk1.pcpi_mul_rs2 [23]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_487 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49234 (.A0
       (\genblk1.pcpi_mul_rs1 [22]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_170 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_95 ), .B1
       (\genblk1.pcpi_mul_rs2 [5]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_486 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49235 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_197 ), .A1
       (\genblk1.pcpi_mul_rs1 [16]), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_89 ), .B1
       (\genblk1.pcpi_mul_rs2 [29]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_485 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49236 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_164 ), .A1
       (\genblk1.pcpi_mul_rs1 [3]), .B0 (\genblk1.pcpi_mul_rs2 [19]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_93 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_484 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49237 (.A0
       (\genblk1.pcpi_mul_rs1 [31]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_43 ), .B1
       (\genblk1.pcpi_mul_rs2 [11]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_483 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49238 (.A0
       (\genblk1.pcpi_mul_rs1 [17]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_83 ), .B1
       (\genblk1.pcpi_mul_rs2 [23]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_482 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49239 (.A0
       (\genblk1.pcpi_mul_rs1 [22]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_95 ), .B1
       (\genblk1.pcpi_mul_rs2 [23]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_481 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49240 (.A0
       (\genblk1.pcpi_mul_rs1 [17]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_163 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_83 ), .B1
       (\genblk1.pcpi_mul_rs2 [9]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_480 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49241 (.A0
       (\genblk1.pcpi_mul_rs1 [20]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_165 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_87 ), .B1
       (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_479 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49242 (.A0
       (\genblk1.pcpi_mul_rs1 [25]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_167 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_53 ), .B1
       (\genblk1.pcpi_mul_rs2 [7]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_478 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49243 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_197 ), .A1
       (\genblk1.pcpi_mul_rs1 [11]), .B0 (\genblk1.pcpi_mul_rs2 [29]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_51 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_477 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49244 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_197 ), .A1
       (\genblk1.pcpi_mul_rs1 [17]), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_83 ), .B1
       (\genblk1.pcpi_mul_rs2 [29]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_476 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49245 (.A0
       (\genblk1.pcpi_mul_rs1 [14]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_163 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_39 ), .B1
       (\genblk1.pcpi_mul_rs2 [9]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_475 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49246 (.A0
       (\genblk1.pcpi_mul_rs1 [29]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_197 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_61 ), .B1
       (\genblk1.pcpi_mul_rs2 [29]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_474 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49247 (.A0
       (\genblk1.pcpi_mul_rs1 [31]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_164 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_43 ), .B1
       (\genblk1.pcpi_mul_rs2 [19]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_473 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49248 (.A0
       (\genblk1.pcpi_mul_rs1 [8]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_196 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_85 ), .B1
       (\genblk1.pcpi_mul_rs2 [13]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_472 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49249 (.A0
       (\genblk1.pcpi_mul_rs1 [29]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_61 ), .B1
       (\genblk1.pcpi_mul_rs2 [23]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_471 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49250 (.A0
       (\genblk1.pcpi_mul_rs1 [11]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_196 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_51 ), .B1
       (\genblk1.pcpi_mul_rs2 [13]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_470 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49251 (.A0
       (\genblk1.pcpi_mul_rs1 [5]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_166 ), .B0
       (\genblk1.pcpi_mul_rs2 [15]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_47 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_469 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49252 (.A0
       (\genblk1.pcpi_mul_rs1 [3]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_196 ), .B0
       (\genblk1.pcpi_mul_rs2 [13]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_93 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_468 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49253 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ), .A1
       (\genblk1.pcpi_mul_rs1 [11]), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_51 ), .B1
       (\genblk1.pcpi_mul_rs2 [23]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_467 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49254 (.A0
       (\genblk1.pcpi_mul_rs1 [24]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_99 ), .B1
       (\genblk1.pcpi_mul_rs2 [11]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_466 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49255 (.A0
       (\genblk1.pcpi_mul_rs1 [26]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_55 ), .B1
       (\genblk1.pcpi_mul_rs2 [11]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_465 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49256 (.A0
       (\genblk1.pcpi_mul_rs1 [30]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_63 ), .B1
       (\genblk1.pcpi_mul_rs2 [11]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_464 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49257 (.A0
       (\genblk1.pcpi_mul_rs1 [14]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_167 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_39 ), .B1
       (\genblk1.pcpi_mul_rs2 [7]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_463 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49258 (.A0
       (\genblk1.pcpi_mul_rs1 [15]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_170 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_97 ), .B1
       (\genblk1.pcpi_mul_rs2 [5]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_462 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49259 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_197 ), .A1
       (\genblk1.pcpi_mul_rs1 [6]), .B0 (\genblk1.pcpi_mul_rs2 [29]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_59 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_461 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49260 (.A0
       (\genblk1.pcpi_mul_rs1 [28]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_197 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_65 ), .B1
       (\genblk1.pcpi_mul_rs2 [29]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_460 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49261 (.A0
       (\genblk1.pcpi_mul_rs1 [29]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_170 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_61 ), .B1
       (\genblk1.pcpi_mul_rs2 [5]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_459 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49262 (.A0
       (\genblk1.pcpi_mul_rs1 [2]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ), .B0
       (\genblk1.pcpi_mul_rs2 [11]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_57 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_458 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49263 (.A0
       (\genblk1.pcpi_mul_rs1 [27]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_77 ), .B1
       (\genblk1.pcpi_mul_rs2 [23]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_457 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49264 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ), .A1
       (\genblk1.pcpi_mul_rs1 [2]), .B0 (\genblk1.pcpi_mul_rs2 [23]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_57 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_456 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49265 (.A0
       (\genblk1.pcpi_mul_rs1 [30]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_167 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_63 ), .B1
       (\genblk1.pcpi_mul_rs2 [7]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_455 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49266 (.A0
       (\genblk1.pcpi_mul_rs1 [15]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_167 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_97 ), .B1
       (\genblk1.pcpi_mul_rs2 [7]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_454 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49267 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_166 ), .A1
       (\genblk1.pcpi_mul_rs1 [1]), .B0 (\genblk1.pcpi_mul_rs2 [15]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_81 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_453 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49268 (.A0
       (\genblk1.pcpi_mul_rs1 [23]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_163 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_49 ), .B1
       (\genblk1.pcpi_mul_rs2 [9]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_452 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49269 (.A0
       (\genblk1.pcpi_mul_rs1 [12]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_167 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_45 ), .B1
       (\genblk1.pcpi_mul_rs2 [7]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_451 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49270 (.A0
       (\genblk1.pcpi_mul_rs1 [13]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_166 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_41 ), .B1
       (\genblk1.pcpi_mul_rs2 [15]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_450 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49271 (.A0
       (\genblk1.pcpi_mul_rs1 [9]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_165 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_75 ), .B1
       (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_449 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49272 (.A0
       (\genblk1.pcpi_mul_rs1 [21]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_195 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_67 ), .B1
       (\genblk1.pcpi_mul_rs2 [21]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_448 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49273 (.A0
       (\genblk1.pcpi_mul_rs1 [7]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_91 ), .B1
       (\genblk1.pcpi_mul_rs2 [11]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_447 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49274 (.A0
       (\genblk1.pcpi_mul_rs1 [22]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_167 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_95 ), .B1
       (\genblk1.pcpi_mul_rs2 [7]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_446 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49275 (.A0
       (\genblk1.pcpi_mul_rs1 [5]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_165 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_47 ), .B1
       (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_445 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49276 (.A0
       (\genblk1.pcpi_mul_rs1 [9]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_163 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_75 ), .B1
       (\genblk1.pcpi_mul_rs2 [9]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_444 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49277 (.A0
       (\genblk1.pcpi_mul_rs1 [21]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_67 ), .B1
       (\genblk1.pcpi_mul_rs2 [23]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_443 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49278 (.A0
       (\genblk1.pcpi_mul_rs1 [29]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_167 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_61 ), .B1
       (\genblk1.pcpi_mul_rs2 [7]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_442 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49279 (.A0
       (\genblk1.pcpi_mul_rs1 [26]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_167 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_55 ), .B1
       (\genblk1.pcpi_mul_rs2 [7]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_441 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49280 (.A0
       (\genblk1.pcpi_mul_rs1 [31]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_166 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_43 ), .B1
       (\genblk1.pcpi_mul_rs2 [15]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_440 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49281 (.A0
       (\genblk1.pcpi_mul_rs1 [1]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ), .B0
       (\genblk1.pcpi_mul_rs2 [11]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_81 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_439 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49282 (.A0
       (\genblk1.pcpi_mul_rs1 [10]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_164 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_69 ), .B1
       (\genblk1.pcpi_mul_rs2 [19]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_438 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49283 (.A0
       (\genblk1.pcpi_mul_rs1 [27]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_193 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_77 ), .B1
       (\genblk1.pcpi_mul_rs2 [27]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_437 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49284 (.A0
       (\genblk1.pcpi_mul_rs1 [8]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_194 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_85 ), .B1
       (\genblk1.pcpi_mul_rs2 [17]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_436 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49285 (.A0
       (\genblk1.pcpi_mul_rs1 [20]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_87 ), .B1
       (\genblk1.pcpi_mul_rs2 [11]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_435 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49286 (.A0
       (\genblk1.pcpi_mul_rs1 [7]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_163 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_91 ), .B1
       (\genblk1.pcpi_mul_rs2 [9]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_434 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49287 (.A0
       (\genblk1.pcpi_mul_rs1 [15]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_163 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_97 ), .B1
       (\genblk1.pcpi_mul_rs2 [9]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_433 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49288 (.A0
       (\genblk1.pcpi_mul_rs1 [3]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_163 ), .B0
       (\genblk1.pcpi_mul_rs2 [9]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_93 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_432 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49289 (.A0
       (\genblk1.pcpi_mul_rs1 [2]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_166 ), .B0
       (\genblk1.pcpi_mul_rs2 [15]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_57 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_431 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49290 (.A0
       (\genblk1.pcpi_mul_rs1 [7]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_170 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_91 ), .B1
       (\genblk1.pcpi_mul_rs2 [5]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_430 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49291 (.A0
       (\genblk1.pcpi_mul_rs1 [20]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_170 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_87 ), .B1
       (\genblk1.pcpi_mul_rs2 [5]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_429 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49292 (.A0
       (\genblk1.pcpi_mul_rs1 [15]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_194 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_97 ), .B1
       (\genblk1.pcpi_mul_rs2 [17]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_428 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49293 (.A0
       (\genblk1.pcpi_mul_rs1 [30]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_163 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_63 ), .B1
       (\genblk1.pcpi_mul_rs2 [9]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_427 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49294 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_197 ), .A1
       (\genblk1.pcpi_mul_rs1 [2]), .B0 (\genblk1.pcpi_mul_rs2 [29]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_57 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_426 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49295 (.A0
       (\genblk1.pcpi_mul_rs1 [4]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_165 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_71 ), .B1
       (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_425 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49296 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_198 ), .A1
       (\genblk1.pcpi_mul_rs1 [17]), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_83 ), .B1
       (\genblk1.pcpi_mul_rs2 [25]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_424 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49297 (.A0
       (\genblk1.pcpi_mul_rs1 [4]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_196 ), .B0
       (\genblk1.pcpi_mul_rs2 [13]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_71 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_423 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49298 (.A0
       (\genblk1.pcpi_mul_rs1 [19]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_194 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_73 ), .B1
       (\genblk1.pcpi_mul_rs2 [17]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_422 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49299 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_198 ), .A1
       (\genblk1.pcpi_mul_rs1 [13]), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_41 ), .B1
       (\genblk1.pcpi_mul_rs2 [25]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_421 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49300 (.A0
       (\genblk1.pcpi_mul_rs1 [17]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_194 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_83 ), .B1
       (\genblk1.pcpi_mul_rs2 [17]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_420 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49301 (.A0
       (\genblk1.pcpi_mul_rs1 [10]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_166 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_69 ), .B1
       (\genblk1.pcpi_mul_rs2 [15]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_419 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49302 (.A0
       (\genblk1.pcpi_mul_rs1 [14]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_170 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_39 ), .B1
       (\genblk1.pcpi_mul_rs2 [5]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_418 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49303 (.A0
       (\genblk1.pcpi_mul_rs1 [14]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_165 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_39 ), .B1
       (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_417 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49304 (.A0
       (\genblk1.pcpi_mul_rs1 [12]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_164 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_45 ), .B1
       (\genblk1.pcpi_mul_rs2 [19]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_416 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49305 (.A0
       (\genblk1.pcpi_mul_rs1 [30]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_196 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_63 ), .B1
       (\genblk1.pcpi_mul_rs2 [13]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_415 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49306 (.A0
       (\genblk1.pcpi_mul_rs1 [21]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_197 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_67 ), .B1
       (\genblk1.pcpi_mul_rs2 [29]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_414 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49307 (.A0
       (\genblk1.pcpi_mul_rs1 [21]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_198 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_67 ), .B1
       (\genblk1.pcpi_mul_rs2 [25]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_413 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49308 (.A0
       (\genblk1.pcpi_mul_rs1 [29]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_163 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_61 ), .B1
       (\genblk1.pcpi_mul_rs2 [9]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_412 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49309 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_198 ), .A1
       (\genblk1.pcpi_mul_rs1 [11]), .B0 (\genblk1.pcpi_mul_rs2 [25]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_51 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_411 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49310 (.A0
       (\genblk1.pcpi_mul_rs1 [19]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_170 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_73 ), .B1
       (\genblk1.pcpi_mul_rs2 [5]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_410 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49311 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_198 ), .A1
       (\genblk1.pcpi_mul_rs1 [18]), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_79 ), .B1
       (\genblk1.pcpi_mul_rs2 [25]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_409 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49312 (.A0
       (\genblk1.pcpi_mul_rs1 [5]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_167 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_47 ), .B1
       (\genblk1.pcpi_mul_rs2 [7]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_408 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49313 (.A0
       (\genblk1.pcpi_mul_rs1 [14]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_194 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_39 ), .B1
       (\genblk1.pcpi_mul_rs2 [17]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_407 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49314 (.A0
       (\genblk1.pcpi_mul_rs1 [18]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_170 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_79 ), .B1
       (\genblk1.pcpi_mul_rs2 [5]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_406 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49315 (.A0
       (\genblk1.pcpi_mul_rs1 [1]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_163 ), .B0
       (\genblk1.pcpi_mul_rs2 [9]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_81 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_405 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49316 (.A0
       (\genblk1.pcpi_mul_rs1 [12]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_170 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_45 ), .B1
       (\genblk1.pcpi_mul_rs2 [5]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_404 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49317 (.A0
       (\genblk1.pcpi_mul_rs1 [7]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_165 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_91 ), .B1
       (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_403 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49318 (.A0
       (\genblk1.pcpi_mul_rs1 [14]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_164 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_39 ), .B1
       (\genblk1.pcpi_mul_rs2 [19]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_402 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49319 (.A0
       (\genblk1.pcpi_mul_rs1 [28]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_167 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_65 ), .B1
       (\genblk1.pcpi_mul_rs2 [7]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_401 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49320 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_198 ), .A1
       (\genblk1.pcpi_mul_rs1 [8]), .B0 (\genblk1.pcpi_mul_rs2 [25]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_85 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_400 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49321 (.A0
       (\genblk1.pcpi_mul_rs1 [8]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_167 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_85 ), .B1
       (\genblk1.pcpi_mul_rs2 [7]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_399 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49322 (.A0
       (\genblk1.pcpi_mul_rs1 [31]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_167 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_43 ), .B1
       (\genblk1.pcpi_mul_rs2 [7]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_398 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49323 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_198 ), .A1
       (\genblk1.pcpi_mul_rs1 [15]), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_97 ), .B1
       (\genblk1.pcpi_mul_rs2 [25]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_397 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49324 (.A0
       (\genblk1.pcpi_mul_rs1 [30]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_193 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_63 ), .B1
       (\genblk1.pcpi_mul_rs2 [27]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_396 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49325 (.A0
       (\genblk1.pcpi_mul_rs1 [20]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_163 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_87 ), .B1
       (\genblk1.pcpi_mul_rs2 [9]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_395 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49326 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_194 ), .A1
       (\genblk1.pcpi_mul_rs1 [2]), .B0 (\genblk1.pcpi_mul_rs2 [17]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_57 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_394 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49327 (.A0
       (\genblk1.pcpi_mul_rs1 [20]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_166 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_87 ), .B1
       (\genblk1.pcpi_mul_rs2 [15]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_393 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49328 (.A0
       (\genblk1.pcpi_mul_rs1 [15]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_195 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_97 ), .B1
       (\genblk1.pcpi_mul_rs2 [21]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_392 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49329 (.A0
       (\genblk1.pcpi_mul_rs1 [31]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_195 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_43 ), .B1
       (\genblk1.pcpi_mul_rs2 [21]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_391 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49330 (.A0
       (\genblk1.pcpi_mul_rs1 [27]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_198 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_77 ), .B1
       (\genblk1.pcpi_mul_rs2 [25]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_390 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49331 (.A0
       (\genblk1.pcpi_mul_rs1 [4]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_163 ), .B0
       (\genblk1.pcpi_mul_rs2 [9]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_71 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_389 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49332 (.A0
       (\genblk1.pcpi_mul_rs1 [24]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_193 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_99 ), .B1
       (\genblk1.pcpi_mul_rs2 [27]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_388 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49333 (.A0
       (\genblk1.pcpi_mul_rs1 [6]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_196 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_59 ), .B1
       (\genblk1.pcpi_mul_rs2 [13]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_387 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49334 (.A0
       (\genblk1.pcpi_mul_rs1 [19]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_164 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_73 ), .B1
       (\genblk1.pcpi_mul_rs2 [19]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_386 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49335 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_197 ), .A1
       (\genblk1.pcpi_mul_rs1 [13]), .B0 (\genblk1.pcpi_mul_rs2 [29]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_41 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_385 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49336 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ), .A1
       (\genblk1.pcpi_mul_rs1 [5]), .B0 (\genblk1.pcpi_mul_rs2 [23]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_47 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_384 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49337 (.A0
       (\genblk1.pcpi_mul_rs1 [20]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_194 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_87 ), .B1
       (\genblk1.pcpi_mul_rs2 [17]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_383 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49338 (.A0
       (\genblk1.pcpi_mul_rs1 [30]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_164 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_63 ), .B1
       (\genblk1.pcpi_mul_rs2 [19]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_382 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49339 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ), .A1
       (\genblk1.pcpi_mul_rs1 [13]), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_41 ), .B1
       (\genblk1.pcpi_mul_rs2 [23]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_381 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49340 (.A0
       (\genblk1.pcpi_mul_rs1 [26]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_197 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_55 ), .B1
       (\genblk1.pcpi_mul_rs2 [29]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_380 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49341 (.A0
       (\genblk1.pcpi_mul_rs1 [3]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_167 ), .B0
       (\genblk1.pcpi_mul_rs2 [7]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_93 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_379 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49342 (.A0
       (\genblk1.pcpi_mul_rs1 [25]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_53 ), .B1
       (\genblk1.pcpi_mul_rs2 [23]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_378 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49343 (.A0
       (\genblk1.pcpi_mul_rs1 [2]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_196 ), .B0
       (\genblk1.pcpi_mul_rs2 [13]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_57 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_377 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49344 (.A0
       (\genblk1.pcpi_mul_rs1 [22]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_194 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_95 ), .B1
       (\genblk1.pcpi_mul_rs2 [17]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_376 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49345 (.A0
       (\genblk1.pcpi_mul_rs1 [7]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_167 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_91 ), .B1
       (\genblk1.pcpi_mul_rs2 [7]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_375 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49346 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ), .A1
       (\genblk1.pcpi_mul_rs1 [14]), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_39 ), .B1
       (\genblk1.pcpi_mul_rs2 [23]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_374 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49347 (.A0
       (\genblk1.pcpi_mul_rs1 [25]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_163 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_53 ), .B1
       (\genblk1.pcpi_mul_rs2 [9]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_373 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49348 (.A0
       (\genblk1.pcpi_mul_rs1 [16]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_167 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_89 ), .B1
       (\genblk1.pcpi_mul_rs2 [7]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_372 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49349 (.A0
       (\genblk1.pcpi_mul_rs1 [11]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_167 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_51 ), .B1
       (\genblk1.pcpi_mul_rs2 [7]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_371 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49350 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ), .A1
       (\genblk1.pcpi_mul_rs1 [12]), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_45 ), .B1
       (\genblk1.pcpi_mul_rs2 [23]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_370 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49351 (.A0
       (\genblk1.pcpi_mul_rs1 [8]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_163 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_85 ), .B1
       (\genblk1.pcpi_mul_rs2 [9]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_369 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49352 (.A0
       (\genblk1.pcpi_mul_rs1 [6]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_163 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_59 ), .B1
       (\genblk1.pcpi_mul_rs2 [9]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_368 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49353 (.A0
       (\genblk1.pcpi_mul_rs1 [25]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_193 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_53 ), .B1
       (\genblk1.pcpi_mul_rs2 [27]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_367 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49354 (.A0
       (\genblk1.pcpi_mul_rs1 [25]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_194 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_53 ), .B1
       (\genblk1.pcpi_mul_rs2 [17]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_366 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49355 (.A0
       (\genblk1.pcpi_mul_rs1 [31]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_170 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_43 ), .B1
       (\genblk1.pcpi_mul_rs2 [5]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_365 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49356 (.A0
       (\genblk1.pcpi_mul_rs1 [8]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_85 ), .B1
       (\genblk1.pcpi_mul_rs2 [11]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_364 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49357 (.A0
       (\genblk1.pcpi_mul_rs1 [26]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_166 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_55 ), .B1
       (\genblk1.pcpi_mul_rs2 [15]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_363 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49358 (.A0
       (\genblk1.pcpi_mul_rs1 [12]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_194 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_45 ), .B1
       (\genblk1.pcpi_mul_rs2 [17]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_362 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49359 (.A0
       (\genblk1.pcpi_mul_rs1 [10]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_170 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_69 ), .B1
       (\genblk1.pcpi_mul_rs2 [5]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_361 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49360 (.A0
       (\genblk1.pcpi_mul_rs1 [22]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_196 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_95 ), .B1
       (\genblk1.pcpi_mul_rs2 [13]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_360 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49361 (.A0
       (\genblk1.pcpi_mul_rs1 [27]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_163 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_77 ), .B1
       (\genblk1.pcpi_mul_rs2 [9]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_359 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49362 (.A0
       (\genblk1.pcpi_mul_rs1 [23]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_49 ), .B1
       (\genblk1.pcpi_mul_rs2 [11]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_358 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49363 (.A0
       (\genblk1.pcpi_mul_rs1 [10]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_165 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_69 ), .B1
       (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_357 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49364 (.A0
       (\genblk1.pcpi_mul_rs1 [19]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_73 ), .B1
       (\genblk1.pcpi_mul_rs2 [23]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_356 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49365 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_193 ), .A1
       (\genblk1.pcpi_mul_rs1 [1]), .B0 (\genblk1.pcpi_mul_rs2 [27]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_81 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_355 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49366 (.A0
       (\genblk1.pcpi_mul_rs1 [22]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_166 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_95 ), .B1
       (\genblk1.pcpi_mul_rs2 [15]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_354 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49367 (.A0
       (\genblk1.pcpi_mul_rs1 [19]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_166 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_73 ), .B1
       (\genblk1.pcpi_mul_rs2 [15]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_353 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49368 (.A0
       (\genblk1.pcpi_mul_rs1 [5]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_47 ), .B1
       (\genblk1.pcpi_mul_rs2 [11]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_352 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49369 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_195 ), .A1
       (\genblk1.pcpi_mul_rs1 [3]), .B0 (\genblk1.pcpi_mul_rs2 [21]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_93 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_351 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49370 (.A0
       (\genblk1.pcpi_mul_rs1 [13]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_167 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_41 ), .B1
       (\genblk1.pcpi_mul_rs2 [7]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_350 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49371 (.A0
       (\genblk1.pcpi_mul_rs1 [24]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_196 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_99 ), .B1
       (\genblk1.pcpi_mul_rs2 [13]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_349 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49372 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .A1
       (\genblk1.pcpi_mul_rs1 [7]), .B0 (\genblk1.pcpi_mul_rs2 [31]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_91 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_348 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49373 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .A1
       (\genblk1.pcpi_mul_rs1 [17]), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_83 ), .B1
       (\genblk1.pcpi_mul_rs2 [31]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_347 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49374 (.A0
       (\genblk1.pcpi_mul_rs1 [6]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_171 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_59 ), .B1
       (\genblk1.pcpi_mul_rs2 [1]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_345 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49375 (.A0
       (\genblk1.pcpi_mul_rs1 [24]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_99 ), .B1
       (\genblk1.pcpi_mul_rs2 [31]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_344 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49376 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .A1
       (\genblk1.pcpi_mul_rs1 [6]), .B0 (\genblk1.pcpi_mul_rs2 [31]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_59 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_343 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49377 (.A0
       (\genblk1.pcpi_mul_rs1 [18]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_171 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_79 ), .B1
       (\genblk1.pcpi_mul_rs2 [1]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_341 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49378 (.A0
       (\genblk1.pcpi_mul_rs1 [8]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_171 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_85 ), .B1
       (\genblk1.pcpi_mul_rs2 [1]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_340 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g49379 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_47 ), .A1
       (\genblk1.pcpi_mul_rs2 [1]), .B0 (\genblk1.pcpi_mul_rs1 [5]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_171 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_338 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49380 (.A0
       (\genblk1.pcpi_mul_rs1 [26]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_171 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_55 ), .B1
       (\genblk1.pcpi_mul_rs2 [1]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_337 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49381 (.A0
       (\genblk1.pcpi_mul_rs1 [9]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_171 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_75 ), .B1
       (\genblk1.pcpi_mul_rs2 [1]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_336 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g49382 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_93 ), .A1
       (\genblk1.pcpi_mul_rs2 [1]), .B0 (\genblk1.pcpi_mul_rs1 [3]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_171 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_334 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49383 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .A1
       (\genblk1.pcpi_mul_rs1 [2]), .B0 (\genblk1.pcpi_mul_rs2 [31]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_57 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_333 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49384 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .A1
       (\genblk1.pcpi_mul_rs1 [19]), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_73 ), .B1
       (\genblk1.pcpi_mul_rs2 [31]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_332 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49385 (.A0
       (\genblk1.pcpi_mul_rs1 [25]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_53 ), .B1
       (\genblk1.pcpi_mul_rs2 [31]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_331 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49386 (.A0
       (\genblk1.pcpi_mul_rs1 [23]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_49 ), .B1
       (\genblk1.pcpi_mul_rs2 [31]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_330 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49387 (.A0
       (\genblk1.pcpi_mul_rs1 [27]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_77 ), .B1
       (\genblk1.pcpi_mul_rs2 [31]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_329 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49388 (.A0
       (\genblk1.pcpi_mul_rs1 [2]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_171 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_57 ), .B1
       (\genblk1.pcpi_mul_rs2 [1]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_327 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49389 (.A0
       (\genblk1.pcpi_mul_rs1 [27]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_171 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_77 ), .B1
       (\genblk1.pcpi_mul_rs2 [1]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_326 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g49390 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_43 ), .A1
       (\genblk1.pcpi_mul_rs2 [1]), .B0 (\genblk1.pcpi_mul_rs1 [31]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_171 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_324 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49391 (.A0
       (\genblk1.pcpi_mul_rs1 [22]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_95 ), .B1
       (\genblk1.pcpi_mul_rs2 [31]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_323 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49392 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .A1
       (\genblk1.pcpi_mul_rs1 [13]), .B0 (\genblk1.pcpi_mul_rs2 [31]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_41 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_322 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g49393 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_91 ), .A1
       (\genblk1.pcpi_mul_rs2 [1]), .B0 (\genblk1.pcpi_mul_rs1 [7]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_171 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_320 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g49394 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_73 ), .A1
       (\genblk1.pcpi_mul_rs2 [1]), .B0 (\genblk1.pcpi_mul_rs1 [19]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_171 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_318 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49395 (.A0
       (\genblk1.pcpi_mul_rs1 [11]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_171 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_51 ), .B1
       (\genblk1.pcpi_mul_rs2 [1]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_317 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49396 (.A0
       (\genblk1.pcpi_mul_rs1 [25]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_171 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_53 ), .B1
       (\genblk1.pcpi_mul_rs2 [1]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_316 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49397 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .A1
       (\genblk1.pcpi_mul_rs1 [3]), .B0 (\genblk1.pcpi_mul_rs2 [31]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_93 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_315 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49398 (.A0
       (\genblk1.pcpi_mul_rs1 [4]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_171 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_71 ), .B1
       (\genblk1.pcpi_mul_rs2 [1]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_313 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49399 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .A1
       (\genblk1.pcpi_mul_rs1 [5]), .B0 (\genblk1.pcpi_mul_rs2 [31]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_47 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_312 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49400 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .A1
       (\genblk1.pcpi_mul_rs1 [4]), .B0 (\genblk1.pcpi_mul_rs2 [31]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_71 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_311 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49401 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .A1
       (\genblk1.pcpi_mul_rs1 [14]), .B0 (\genblk1.pcpi_mul_rs2 [31]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_39 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_310 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49402 (.A0
       (\genblk1.pcpi_mul_rs1 [28]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_65 ), .B1
       (\genblk1.pcpi_mul_rs2 [31]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_309 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49403 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .A1
       (\genblk1.pcpi_mul_rs1 [10]), .B0 (\genblk1.pcpi_mul_rs2 [31]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_69 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_308 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49404 (.A0
       (\genblk1.pcpi_mul_rs1 [31]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_43 ), .B1
       (\genblk1.pcpi_mul_rs2 [31]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_307 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g49405 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_41 ), .A1
       (\genblk1.pcpi_mul_rs2 [1]), .B0 (\genblk1.pcpi_mul_rs1 [13]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_171 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_305 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49406 (.A0
       (\genblk1.pcpi_mul_rs1 [21]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_67 ), .B1
       (\genblk1.pcpi_mul_rs2 [31]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_304 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49407 (.A0
       (\genblk1.pcpi_mul_rs1 [20]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_171 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_87 ), .B1
       (\genblk1.pcpi_mul_rs2 [1]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_303 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49408 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .A1
       (\genblk1.pcpi_mul_rs1 [8]), .B0 (\genblk1.pcpi_mul_rs2 [31]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_85 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_302 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49409 (.A0
       (\genblk1.pcpi_mul_rs1 [21]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_171 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_67 ), .B1
       (\genblk1.pcpi_mul_rs2 [1]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_301 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49410 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .A1
       (\genblk1.pcpi_mul_rs1 [12]), .B0 (\genblk1.pcpi_mul_rs2 [31]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_45 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_300 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g49411 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_83 ), .A1
       (\genblk1.pcpi_mul_rs2 [1]), .B0 (\genblk1.pcpi_mul_rs1 [17]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_171 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_298 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49412 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .A1
       (\genblk1.pcpi_mul_rs1 [1]), .B0 (\genblk1.pcpi_mul_rs2 [31]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_81 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_297 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49413 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .A1
       (\genblk1.pcpi_mul_rs1 [11]), .B0 (\genblk1.pcpi_mul_rs2 [31]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_51 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_296 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49414 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .A1
       (\genblk1.pcpi_mul_rs1 [15]), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_97 ), .B1
       (\genblk1.pcpi_mul_rs2 [31]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_295 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49415 (.A0
       (\genblk1.pcpi_mul_rs1 [28]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_171 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_65 ), .B1
       (\genblk1.pcpi_mul_rs2 [1]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_293 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49416 (.A0
       (\genblk1.pcpi_mul_rs1 [30]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_63 ), .B1
       (\genblk1.pcpi_mul_rs2 [31]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_292 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49417 (.A0
       (\genblk1.pcpi_mul_rs1 [24]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_171 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_99 ), .B1
       (\genblk1.pcpi_mul_rs2 [1]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_291 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g49418 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_63 ), .A1
       (\genblk1.pcpi_mul_rs2 [1]), .B0 (\genblk1.pcpi_mul_rs1 [30]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_171 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_289 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49419 (.A0
       (\genblk1.pcpi_mul_rs1 [26]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_55 ), .B1
       (\genblk1.pcpi_mul_rs2 [31]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_288 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49420 (.A0
       (\genblk1.pcpi_mul_rs1 [14]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_171 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_39 ), .B1
       (\genblk1.pcpi_mul_rs2 [1]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_286 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49421 (.A0
       (\genblk1.pcpi_mul_rs1 [10]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_171 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_69 ), .B1
       (\genblk1.pcpi_mul_rs2 [1]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_285 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49422 (.A0
       (\genblk1.pcpi_mul_rs1 [23]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_171 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_49 ), .B1
       (\genblk1.pcpi_mul_rs2 [1]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_284 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49423 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .A1
       (\genblk1.pcpi_mul_rs1 [16]), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_89 ), .B1
       (\genblk1.pcpi_mul_rs2 [31]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_283 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g49424 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_97 ), .A1
       (\genblk1.pcpi_mul_rs2 [1]), .B0 (\genblk1.pcpi_mul_rs1 [15]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_171 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_281 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g49425 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_81 ), .A1
       (\genblk1.pcpi_mul_rs2 [1]), .B0 (\genblk1.pcpi_mul_rs1 [1]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_171 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_279 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49426 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .A1
       (\genblk1.pcpi_mul_rs1 [9]), .B0 (\genblk1.pcpi_mul_rs2 [31]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_75 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_278 ));
  OAI22X1 \genblk1.pcpi_mul_mul_2366_47_g49427 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_61 ), .A1
       (\genblk1.pcpi_mul_rs2 [1]), .B0 (\genblk1.pcpi_mul_rs1 [29]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_171 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_276 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49428 (.A0
       (\genblk1.pcpi_mul_rs1 [20]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_87 ), .B1
       (\genblk1.pcpi_mul_rs2 [31]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_275 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49429 (.A0
       (\genblk1.pcpi_mul_rs1 [16]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_171 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_89 ), .B1
       (\genblk1.pcpi_mul_rs2 [1]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_273 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49430 (.A0
       (\genblk1.pcpi_mul_rs1 [29]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_61 ), .B1
       (\genblk1.pcpi_mul_rs2 [31]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_272 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49431 (.A0
       (\genblk1.pcpi_mul_rs1 [12]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_171 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_45 ), .B1
       (\genblk1.pcpi_mul_rs2 [1]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_270 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49432 (.A0
       (\genblk1.pcpi_mul_rs1 [22]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_171 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_95 ), .B1
       (\genblk1.pcpi_mul_rs2 [1]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_269 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49433 (.A0
       (\genblk1.pcpi_mul_rs1 [18]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_79 ), .B1
       (\genblk1.pcpi_mul_rs2 [31]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_268 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49434 (.A0
       (\genblk1.pcpi_mul_rs1 [28]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_65 ), .B1
       (\genblk1.pcpi_mul_rs2 [11]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_267 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49435 (.A0
       (\genblk1.pcpi_mul_rs1 [4]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_167 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_71 ), .B1
       (\genblk1.pcpi_mul_rs2 [7]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_266 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49436 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_197 ), .A1
       (\genblk1.pcpi_mul_rs1 [3]), .B0 (\genblk1.pcpi_mul_rs2 [29]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_93 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_265 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49437 (.A0
       (\genblk1.pcpi_mul_rs1 [9]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_167 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_75 ), .B1
       (\genblk1.pcpi_mul_rs2 [7]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_264 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49438 (.A0
       (\genblk1.pcpi_mul_rs1 [30]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_195 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_63 ), .B1
       (\genblk1.pcpi_mul_rs2 [21]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_263 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49439 (.A0
       (\genblk1.pcpi_mul_rs1 [28]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_65 ), .B1
       (\genblk1.pcpi_mul_rs2 [23]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_262 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49440 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_198 ), .A1
       (\genblk1.pcpi_mul_rs1 [12]), .B0 (\genblk1.pcpi_mul_rs2 [25]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_45 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_261 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49441 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_193 ), .A1
       (\genblk1.pcpi_mul_rs1 [3]), .B0 (\genblk1.pcpi_mul_rs2 [27]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_93 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_260 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49442 (.A0
       (\genblk1.pcpi_mul_rs1 [16]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_170 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_89 ), .B1
       (\genblk1.pcpi_mul_rs2 [5]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_259 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49443 (.A0
       (\genblk1.pcpi_mul_rs1 [9]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_166 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_75 ), .B1
       (\genblk1.pcpi_mul_rs2 [15]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_258 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49444 (.A0
       (\genblk1.pcpi_mul_rs1 [2]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_170 ), .B0
       (\genblk1.pcpi_mul_rs2 [5]), .B1
       (\genblk1.pcpi_mul_mul_2366_47_n_57 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_257 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49445 (.A0
       (\genblk1.pcpi_mul_rs1 [18]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_165 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_79 ), .B1
       (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_256 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49446 (.A0
       (\genblk1.pcpi_mul_rs1 [31]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_194 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_43 ), .B1
       (\genblk1.pcpi_mul_rs2 [17]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_255 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49447 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ), .A1
       (\genblk1.pcpi_mul_rs1 [1]), .B0 (\genblk1.pcpi_mul_rs2 [23]),
       .B1 (\genblk1.pcpi_mul_mul_2366_47_n_81 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_254 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49448 (.A0
       (\genblk1.pcpi_mul_rs1 [24]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_198 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_99 ), .B1
       (\genblk1.pcpi_mul_rs2 [25]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_253 ));
  AOI22X1 \genblk1.pcpi_mul_mul_2366_47_g49449 (.A0
       (\genblk1.pcpi_mul_rs1 [13]), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_41 ), .B1
       (\genblk1.pcpi_mul_rs2 [11]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_252 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_g49457 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_224 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_223 ));
  NOR2X1 \genblk1.pcpi_mul_mul_2366_47_g49458 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_37 ), .B
       (\genblk1.pcpi_mul_rs2 [1]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_228 ));
  NAND2X1 \genblk1.pcpi_mul_mul_2366_47_g49460 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_172 ), .B
       (\genblk1.pcpi_mul_rs2 [31]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_221 ));
  NOR2X1 \genblk1.pcpi_mul_mul_2366_47_g49461 (.A
       (\genblk1.pcpi_mul_rs1 [32]), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_171 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_227 ));
  NAND2X1 \genblk1.pcpi_mul_mul_2366_47_g49463 (.A
       (\genblk1.pcpi_mul_rs2 [32]), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_226 ));
  NOR2X1 \genblk1.pcpi_mul_mul_2366_47_g49464 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_35 ), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .Y
       (\genblk1.pcpi_mul_n_91 ));
  OR2X1 \genblk1.pcpi_mul_mul_2366_47_g49465 (.A
       (\genblk1.pcpi_mul_rs2 [0]), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_171 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_224 ));
  INVX2 \genblk1.pcpi_mul_mul_2366_47_g49491 (.A
       (\genblk1.pcpi_mul_rs2 [31]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_199 ));
  INVX2 \genblk1.pcpi_mul_mul_2366_47_g49492 (.A
       (\genblk1.pcpi_mul_rs2 [25]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_198 ));
  INVX2 \genblk1.pcpi_mul_mul_2366_47_g49493 (.A
       (\genblk1.pcpi_mul_rs2 [29]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_197 ));
  INVX2 \genblk1.pcpi_mul_mul_2366_47_g49494 (.A
       (\genblk1.pcpi_mul_rs2 [13]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_196 ));
  INVX2 \genblk1.pcpi_mul_mul_2366_47_g49495 (.A
       (\genblk1.pcpi_mul_rs2 [21]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_195 ));
  INVX2 \genblk1.pcpi_mul_mul_2366_47_g49496 (.A
       (\genblk1.pcpi_mul_rs2 [17]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_194 ));
  INVX2 \genblk1.pcpi_mul_mul_2366_47_g49497 (.A
       (\genblk1.pcpi_mul_rs2 [27]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_193 ));
  INVX2 \genblk1.pcpi_mul_mul_2366_47_g49523 (.A
       (\genblk1.pcpi_mul_rs2 [1]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_171 ));
  INVX2 \genblk1.pcpi_mul_mul_2366_47_g49524 (.A
       (\genblk1.pcpi_mul_rs2 [5]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_170 ));
  INVX2 \genblk1.pcpi_mul_mul_2366_47_g49525 (.A
       (\genblk1.pcpi_mul_rs2 [11]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_169 ));
  INVX2 \genblk1.pcpi_mul_mul_2366_47_g49526 (.A
       (\genblk1.pcpi_mul_rs2 [23]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_168 ));
  INVX2 \genblk1.pcpi_mul_mul_2366_47_g49527 (.A
       (\genblk1.pcpi_mul_rs2 [7]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_167 ));
  INVX2 \genblk1.pcpi_mul_mul_2366_47_g49528 (.A
       (\genblk1.pcpi_mul_rs2 [15]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_166 ));
  INVX2 \genblk1.pcpi_mul_mul_2366_47_g49529 (.A
       (\genblk1.pcpi_mul_rs2 [3]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_165 ));
  INVX2 \genblk1.pcpi_mul_mul_2366_47_g49530 (.A
       (\genblk1.pcpi_mul_rs2 [19]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_164 ));
  INVX2 \genblk1.pcpi_mul_mul_2366_47_g49531 (.A
       (\genblk1.pcpi_mul_rs2 [9]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_163 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_drc_bufs49538 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_569 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_156 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_drc_bufs49545 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_157 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_drc_bufs49552 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_150 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_drc_bufs49559 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_148 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_drc_bufs49566 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_147 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_drc_bufs49573 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_161 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_drc_bufs49580 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_160 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_drc_bufs49587 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_149 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_drc_bufs49594 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_159 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_drc_bufs49601 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_151 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_drc_bufs49608 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_158 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_drc_bufs49615 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_155 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_drc_bufs49622 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_153 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_drc_bufs49629 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_152 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_drc_bufs49636 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_154 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_drc_bufs49748 (.A
       (\genblk1.pcpi_mul_mul_2366_47_n_137 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_162 ));
  INVX3 \genblk1.pcpi_mul_mul_2366_47_drc_bufs49874 (.A
       (\genblk1.pcpi_mul_rs1 [0]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_drc_bufs50142 (.A
       (\genblk1.pcpi_mul_rs2 [10]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_24 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_drc_bufs50146 (.A
       (\genblk1.pcpi_mul_rs2 [26]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_22 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_drc_bufs50150 (.A
       (\genblk1.pcpi_mul_rs2 [20]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_20 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_drc_bufs50154 (.A
       (\genblk1.pcpi_mul_rs2 [22]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_18 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_drc_bufs50158 (.A
       (\genblk1.pcpi_mul_rs2 [24]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_16 ));
  INVX1 \genblk1.pcpi_mul_mul_2366_47_drc_bufs50162 (.A
       (\genblk1.pcpi_mul_rs2 [8]), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_14 ));
  AO21X1 \genblk1.pcpi_mul_mul_2366_47_g2 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_563 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_827 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_803 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_13 ));
  AO21X1 \genblk1.pcpi_mul_mul_2366_47_g50164 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_574 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_826 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_802 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_12 ));
  AO21X1 \genblk1.pcpi_mul_mul_2366_47_g50165 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_565 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_830 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_801 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_11 ));
  AO21X1 \genblk1.pcpi_mul_mul_2366_47_g50166 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_564 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_829 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_800 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_10 ));
  AO21X1 \genblk1.pcpi_mul_mul_2366_47_g50167 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_573 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_831 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_799 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_9 ));
  AO21X1 \genblk1.pcpi_mul_mul_2366_47_g50168 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_570 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_833 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_798 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_8 ));
  AO21X1 \genblk1.pcpi_mul_mul_2366_47_g50169 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_568 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_832 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_797 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_7 ));
  AO21X1 \genblk1.pcpi_mul_mul_2366_47_g50170 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_562 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_824 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_796 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_6 ));
  AO21X1 \genblk1.pcpi_mul_mul_2366_47_g50171 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_567 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_828 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_795 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_5 ));
  AO21X1 \genblk1.pcpi_mul_mul_2366_47_g50172 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_560 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_834 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_794 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_4 ));
  AO21X1 \genblk1.pcpi_mul_mul_2366_47_g50173 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_572 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_823 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_793 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_3 ));
  AO21X1 \genblk1.pcpi_mul_mul_2366_47_g50174 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_571 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_825 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_792 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_2 ));
  AO21X1 \genblk1.pcpi_mul_mul_2366_47_g50175 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_566 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_822 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_791 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_1 ));
  AO21X1 \genblk1.pcpi_mul_mul_2366_47_g50176 (.A0
       (\genblk1.pcpi_mul_mul_2366_47_n_561 ), .A1
       (\genblk1.pcpi_mul_mul_2366_47_n_835 ), .B0
       (\genblk1.pcpi_mul_mul_2366_47_n_790 ), .Y
       (\genblk1.pcpi_mul_mul_2366_47_n_0 ));
  AND2X1 \genblk2.pcpi_div_lte_2493_16_g1379 (.A
       (\genblk2.pcpi_div_lte_2493_16_n_102 ), .B
       (\genblk2.pcpi_div_lte_2493_16_n_65 ), .Y
       (\genblk2.pcpi_div_n_314 ));
  NOR4X1 \genblk2.pcpi_div_lte_2493_16_g1380 (.A
       (\genblk2.pcpi_div_divisor [57]), .B
       (\genblk2.pcpi_div_divisor [56]), .C
       (\genblk2.pcpi_div_divisor [58]), .D
       (\genblk2.pcpi_div_lte_2493_16_n_101 ), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_102 ));
  NAND4XL \genblk2.pcpi_div_lte_2493_16_g1381 (.A
       (\genblk2.pcpi_div_lte_2493_16_n_64 ), .B
       (\genblk2.pcpi_div_lte_2493_16_n_62 ), .C
       (\genblk2.pcpi_div_lte_2493_16_n_66 ), .D
       (\genblk2.pcpi_div_lte_2493_16_n_100 ), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_101 ));
  NOR4X1 \genblk2.pcpi_div_lte_2493_16_g1382 (.A
       (\genblk2.pcpi_div_divisor [40]), .B
       (\genblk2.pcpi_div_divisor [39]), .C
       (\genblk2.pcpi_div_divisor [41]), .D
       (\genblk2.pcpi_div_lte_2493_16_n_99 ), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_100 ));
  NAND2X1 \genblk2.pcpi_div_lte_2493_16_g1383 (.A
       (\genblk2.pcpi_div_lte_2493_16_n_61 ), .B
       (\genblk2.pcpi_div_lte_2493_16_n_98 ), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_99 ));
  NOR4X1 \genblk2.pcpi_div_lte_2493_16_g1384 (.A
       (\genblk2.pcpi_div_divisor [32]), .B
       (\genblk2.pcpi_div_divisor [33]), .C
       (\genblk2.pcpi_div_lte_2493_16_n_53 ), .D
       (\genblk2.pcpi_div_lte_2493_16_n_97 ), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_98 ));
  AOI22X1 \genblk2.pcpi_div_lte_2493_16_g1385 (.A0
       (\genblk2.pcpi_div_lte_2493_16_n_56 ), .A1
       (\genblk2.pcpi_div_lte_2493_16_n_96 ), .B0
       (\genblk2.pcpi_div_lte_2493_16_n_9 ), .B1
       (\genblk2.pcpi_div_dividend [31]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_97 ));
  OAI222X1 \genblk2.pcpi_div_lte_2493_16_g1386 (.A0
       (\genblk2.pcpi_div_divisor [30]), .A1
       (\genblk2.pcpi_div_lte_2493_16_n_29 ), .B0
       (\genblk2.pcpi_div_lte_2493_16_n_49 ), .B1
       (\genblk2.pcpi_div_lte_2493_16_n_95 ), .C0
       (\genblk2.pcpi_div_divisor [29]), .C1
       (\genblk2.pcpi_div_lte_2493_16_n_7 ), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_96 ));
  AOI22X1 \genblk2.pcpi_div_lte_2493_16_g1387 (.A0
       (\genblk2.pcpi_div_lte_2493_16_n_30 ), .A1
       (\genblk2.pcpi_div_lte_2493_16_n_94 ), .B0
       (\genblk2.pcpi_div_lte_2493_16_n_4 ), .B1
       (\genblk2.pcpi_div_dividend [28]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_95 ));
  OAI22X1 \genblk2.pcpi_div_lte_2493_16_g1388 (.A0
       (\genblk2.pcpi_div_lte_2493_16_n_31 ), .A1
       (\genblk2.pcpi_div_lte_2493_16_n_93 ), .B0
       (\genblk2.pcpi_div_divisor [27]), .B1
       (\genblk2.pcpi_div_lte_2493_16_n_21 ), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_94 ));
  AOI22X1 \genblk2.pcpi_div_lte_2493_16_g1389 (.A0
       (\genblk2.pcpi_div_lte_2493_16_n_38 ), .A1
       (\genblk2.pcpi_div_lte_2493_16_n_92 ), .B0
       (\genblk2.pcpi_div_lte_2493_16_n_12 ), .B1
       (\genblk2.pcpi_div_dividend [26]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_93 ));
  OAI22X1 \genblk2.pcpi_div_lte_2493_16_g1390 (.A0
       (\genblk2.pcpi_div_lte_2493_16_n_46 ), .A1
       (\genblk2.pcpi_div_lte_2493_16_n_91 ), .B0
       (\genblk2.pcpi_div_divisor [25]), .B1
       (\genblk2.pcpi_div_lte_2493_16_n_3 ), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_92 ));
  AOI22X1 \genblk2.pcpi_div_lte_2493_16_g1391 (.A0
       (\genblk2.pcpi_div_lte_2493_16_n_34 ), .A1
       (\genblk2.pcpi_div_lte_2493_16_n_90 ), .B0
       (\genblk2.pcpi_div_lte_2493_16_n_25 ), .B1
       (\genblk2.pcpi_div_dividend [24]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_91 ));
  OAI22X1 \genblk2.pcpi_div_lte_2493_16_g1392 (.A0
       (\genblk2.pcpi_div_lte_2493_16_n_50 ), .A1
       (\genblk2.pcpi_div_lte_2493_16_n_89 ), .B0
       (\genblk2.pcpi_div_divisor [23]), .B1
       (\genblk2.pcpi_div_lte_2493_16_n_0 ), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_90 ));
  AOI22X1 \genblk2.pcpi_div_lte_2493_16_g1393 (.A0
       (\genblk2.pcpi_div_lte_2493_16_n_39 ), .A1
       (\genblk2.pcpi_div_lte_2493_16_n_88 ), .B0
       (\genblk2.pcpi_div_lte_2493_16_n_8 ), .B1
       (\genblk2.pcpi_div_dividend [22]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_89 ));
  OAI22X1 \genblk2.pcpi_div_lte_2493_16_g1394 (.A0
       (\genblk2.pcpi_div_lte_2493_16_n_59 ), .A1
       (\genblk2.pcpi_div_lte_2493_16_n_87 ), .B0
       (\genblk2.pcpi_div_divisor [21]), .B1
       (\genblk2.pcpi_div_lte_2493_16_n_20 ), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_88 ));
  AOI22X1 \genblk2.pcpi_div_lte_2493_16_g1395 (.A0
       (\genblk2.pcpi_div_lte_2493_16_n_58 ), .A1
       (\genblk2.pcpi_div_lte_2493_16_n_86 ), .B0
       (\genblk2.pcpi_div_lte_2493_16_n_15 ), .B1
       (\genblk2.pcpi_div_dividend [20]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_87 ));
  OAI22X1 \genblk2.pcpi_div_lte_2493_16_g1396 (.A0
       (\genblk2.pcpi_div_lte_2493_16_n_57 ), .A1
       (\genblk2.pcpi_div_lte_2493_16_n_85 ), .B0
       (\genblk2.pcpi_div_divisor [19]), .B1
       (\genblk2.pcpi_div_lte_2493_16_n_2 ), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_86 ));
  AOI22X1 \genblk2.pcpi_div_lte_2493_16_g1397 (.A0
       (\genblk2.pcpi_div_lte_2493_16_n_54 ), .A1
       (\genblk2.pcpi_div_lte_2493_16_n_84 ), .B0
       (\genblk2.pcpi_div_lte_2493_16_n_19 ), .B1
       (\genblk2.pcpi_div_dividend [18]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_85 ));
  OAI22X1 \genblk2.pcpi_div_lte_2493_16_g1398 (.A0
       (\genblk2.pcpi_div_lte_2493_16_n_52 ), .A1
       (\genblk2.pcpi_div_lte_2493_16_n_83 ), .B0
       (\genblk2.pcpi_div_divisor [17]), .B1
       (\genblk2.pcpi_div_lte_2493_16_n_24 ), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_84 ));
  AOI22X1 \genblk2.pcpi_div_lte_2493_16_g1399 (.A0
       (\genblk2.pcpi_div_lte_2493_16_n_51 ), .A1
       (\genblk2.pcpi_div_lte_2493_16_n_82 ), .B0
       (\genblk2.pcpi_div_lte_2493_16_n_27 ), .B1
       (\genblk2.pcpi_div_dividend [16]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_83 ));
  OAI22X1 \genblk2.pcpi_div_lte_2493_16_g1400 (.A0
       (\genblk2.pcpi_div_lte_2493_16_n_48 ), .A1
       (\genblk2.pcpi_div_lte_2493_16_n_81 ), .B0
       (\genblk2.pcpi_div_divisor [15]), .B1
       (\genblk2.pcpi_div_lte_2493_16_n_5 ), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_82 ));
  AOI22X1 \genblk2.pcpi_div_lte_2493_16_g1401 (.A0
       (\genblk2.pcpi_div_lte_2493_16_n_47 ), .A1
       (\genblk2.pcpi_div_lte_2493_16_n_80 ), .B0
       (\genblk2.pcpi_div_lte_2493_16_n_23 ), .B1
       (\genblk2.pcpi_div_dividend [14]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_81 ));
  OAI22X1 \genblk2.pcpi_div_lte_2493_16_g1402 (.A0
       (\genblk2.pcpi_div_lte_2493_16_n_37 ), .A1
       (\genblk2.pcpi_div_lte_2493_16_n_79 ), .B0
       (\genblk2.pcpi_div_divisor [13]), .B1
       (\genblk2.pcpi_div_lte_2493_16_n_13 ), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_80 ));
  AOI22X1 \genblk2.pcpi_div_lte_2493_16_g1403 (.A0
       (\genblk2.pcpi_div_lte_2493_16_n_43 ), .A1
       (\genblk2.pcpi_div_lte_2493_16_n_78 ), .B0
       (\genblk2.pcpi_div_lte_2493_16_n_16 ), .B1
       (\genblk2.pcpi_div_dividend [12]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_79 ));
  OAI22X1 \genblk2.pcpi_div_lte_2493_16_g1404 (.A0
       (\genblk2.pcpi_div_lte_2493_16_n_32 ), .A1
       (\genblk2.pcpi_div_lte_2493_16_n_77 ), .B0
       (\genblk2.pcpi_div_divisor [11]), .B1
       (\genblk2.pcpi_div_lte_2493_16_n_17 ), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_78 ));
  AOI22X1 \genblk2.pcpi_div_lte_2493_16_g1405 (.A0
       (\genblk2.pcpi_div_lte_2493_16_n_40 ), .A1
       (\genblk2.pcpi_div_lte_2493_16_n_76 ), .B0
       (\genblk2.pcpi_div_lte_2493_16_n_11 ), .B1
       (\genblk2.pcpi_div_dividend [10]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_77 ));
  OAI22X1 \genblk2.pcpi_div_lte_2493_16_g1406 (.A0
       (\genblk2.pcpi_div_lte_2493_16_n_44 ), .A1
       (\genblk2.pcpi_div_lte_2493_16_n_75 ), .B0
       (\genblk2.pcpi_div_divisor [9]), .B1
       (\genblk2.pcpi_div_lte_2493_16_n_6 ), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_76 ));
  AOI22X1 \genblk2.pcpi_div_lte_2493_16_g1407 (.A0
       (\genblk2.pcpi_div_lte_2493_16_n_41 ), .A1
       (\genblk2.pcpi_div_lte_2493_16_n_74 ), .B0
       (\genblk2.pcpi_div_lte_2493_16_n_18 ), .B1
       (\genblk2.pcpi_div_dividend [8]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_75 ));
  OAI22X1 \genblk2.pcpi_div_lte_2493_16_g1408 (.A0
       (\genblk2.pcpi_div_lte_2493_16_n_36 ), .A1
       (\genblk2.pcpi_div_lte_2493_16_n_73 ), .B0
       (\genblk2.pcpi_div_divisor [7]), .B1
       (\genblk2.pcpi_div_lte_2493_16_n_28 ), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_74 ));
  AOI22X1 \genblk2.pcpi_div_lte_2493_16_g1409 (.A0
       (\genblk2.pcpi_div_lte_2493_16_n_60 ), .A1
       (\genblk2.pcpi_div_lte_2493_16_n_72 ), .B0
       (\genblk2.pcpi_div_lte_2493_16_n_26 ), .B1
       (\genblk2.pcpi_div_dividend [6]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_73 ));
  OAI22X1 \genblk2.pcpi_div_lte_2493_16_g1410 (.A0
       (\genblk2.pcpi_div_lte_2493_16_n_33 ), .A1
       (\genblk2.pcpi_div_lte_2493_16_n_71 ), .B0
       (\genblk2.pcpi_div_divisor [5]), .B1
       (\genblk2.pcpi_div_lte_2493_16_n_1 ), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_72 ));
  AOI22X1 \genblk2.pcpi_div_lte_2493_16_g1411 (.A0
       (\genblk2.pcpi_div_lte_2493_16_n_35 ), .A1
       (\genblk2.pcpi_div_lte_2493_16_n_70 ), .B0
       (\genblk2.pcpi_div_lte_2493_16_n_10 ), .B1
       (\genblk2.pcpi_div_dividend [4]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_71 ));
  OAI22X1 \genblk2.pcpi_div_lte_2493_16_g1412 (.A0
       (\genblk2.pcpi_div_lte_2493_16_n_42 ), .A1
       (\genblk2.pcpi_div_lte_2493_16_n_69 ), .B0
       (\genblk2.pcpi_div_divisor [3]), .B1
       (\genblk2.pcpi_div_lte_2493_16_n_14 ), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_70 ));
  AOI22X1 \genblk2.pcpi_div_lte_2493_16_g1413 (.A0
       (\genblk2.pcpi_div_lte_2493_16_n_55 ), .A1
       (\genblk2.pcpi_div_lte_2493_16_n_68 ), .B0
       (\genblk2.pcpi_div_lte_2493_16_n_22 ), .B1
       (\genblk2.pcpi_div_dividend [2]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_69 ));
  OAI21X1 \genblk2.pcpi_div_lte_2493_16_g1414 (.A0
       (\genblk2.pcpi_div_divisor [1]), .A1
       (\genblk2.pcpi_div_lte_2493_16_n_45 ), .B0
       (\genblk2.pcpi_div_lte_2493_16_n_67 ), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_68 ));
  OAI2BB1X1 \genblk2.pcpi_div_lte_2493_16_g1415 (.A0N
       (\genblk2.pcpi_div_divisor [1]), .A1N
       (\genblk2.pcpi_div_lte_2493_16_n_45 ), .B0
       (\genblk2.pcpi_div_dividend [1]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_67 ));
  NOR4X1 \genblk2.pcpi_div_lte_2493_16_g1416 (.A
       (\genblk2.pcpi_div_divisor [38]), .B
       (\genblk2.pcpi_div_divisor [55]), .C
       (\genblk2.pcpi_div_divisor [54]), .D
       (\genblk2.pcpi_div_lte_2493_16_n_63 ), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_66 ));
  NOR4X1 \genblk2.pcpi_div_lte_2493_16_g1417 (.A
       (\genblk2.pcpi_div_divisor [61]), .B
       (\genblk2.pcpi_div_divisor [60]), .C
       (\genblk2.pcpi_div_divisor [62]), .D
       (\genblk2.pcpi_div_divisor [59]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_65 ));
  NOR4X1 \genblk2.pcpi_div_lte_2493_16_g1418 (.A
       (\genblk2.pcpi_div_divisor [48]), .B
       (\genblk2.pcpi_div_divisor [47]), .C
       (\genblk2.pcpi_div_divisor [49]), .D
       (\genblk2.pcpi_div_divisor [46]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_64 ));
  OR4X1 \genblk2.pcpi_div_lte_2493_16_g1419 (.A
       (\genblk2.pcpi_div_divisor [52]), .B
       (\genblk2.pcpi_div_divisor [53]), .C
       (\genblk2.pcpi_div_divisor [50]), .D
       (\genblk2.pcpi_div_divisor [51]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_63 ));
  NOR4X1 \genblk2.pcpi_div_lte_2493_16_g1420 (.A
       (\genblk2.pcpi_div_divisor [44]), .B
       (\genblk2.pcpi_div_divisor [43]), .C
       (\genblk2.pcpi_div_divisor [45]), .D
       (\genblk2.pcpi_div_divisor [42]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_62 ));
  NOR4X1 \genblk2.pcpi_div_lte_2493_16_g1421 (.A
       (\genblk2.pcpi_div_divisor [36]), .B
       (\genblk2.pcpi_div_divisor [35]), .C
       (\genblk2.pcpi_div_divisor [37]), .D
       (\genblk2.pcpi_div_divisor [34]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_61 ));
  NAND2BX1 \genblk2.pcpi_div_lte_2493_16_g1422 (.AN
       (\genblk2.pcpi_div_dividend [6]), .B
       (\genblk2.pcpi_div_divisor [6]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_60 ));
  NOR2BX1 \genblk2.pcpi_div_lte_2493_16_g1423 (.AN
       (\genblk2.pcpi_div_divisor [21]), .B
       (\genblk2.pcpi_div_dividend [21]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_59 ));
  NAND2BX1 \genblk2.pcpi_div_lte_2493_16_g1424 (.AN
       (\genblk2.pcpi_div_dividend [20]), .B
       (\genblk2.pcpi_div_divisor [20]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_58 ));
  NOR2BX1 \genblk2.pcpi_div_lte_2493_16_g1425 (.AN
       (\genblk2.pcpi_div_divisor [19]), .B
       (\genblk2.pcpi_div_dividend [19]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_57 ));
  NAND2X1 \genblk2.pcpi_div_lte_2493_16_g1426 (.A
       (\genblk2.pcpi_div_divisor [30]), .B
       (\genblk2.pcpi_div_lte_2493_16_n_29 ), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_56 ));
  NAND2BX1 \genblk2.pcpi_div_lte_2493_16_g1427 (.AN
       (\genblk2.pcpi_div_dividend [2]), .B
       (\genblk2.pcpi_div_divisor [2]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_55 ));
  NAND2BX1 \genblk2.pcpi_div_lte_2493_16_g1428 (.AN
       (\genblk2.pcpi_div_dividend [18]), .B
       (\genblk2.pcpi_div_divisor [18]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_54 ));
  NOR2X1 \genblk2.pcpi_div_lte_2493_16_g1429 (.A
       (\genblk2.pcpi_div_lte_2493_16_n_9 ), .B
       (\genblk2.pcpi_div_dividend [31]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_53 ));
  NOR2BX1 \genblk2.pcpi_div_lte_2493_16_g1430 (.AN
       (\genblk2.pcpi_div_divisor [17]), .B
       (\genblk2.pcpi_div_dividend [17]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_52 ));
  NAND2BX1 \genblk2.pcpi_div_lte_2493_16_g1431 (.AN
       (\genblk2.pcpi_div_dividend [16]), .B
       (\genblk2.pcpi_div_divisor [16]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_51 ));
  NOR2BX1 \genblk2.pcpi_div_lte_2493_16_g1432 (.AN
       (\genblk2.pcpi_div_divisor [23]), .B
       (\genblk2.pcpi_div_dividend [23]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_50 ));
  NOR2BX1 \genblk2.pcpi_div_lte_2493_16_g1433 (.AN
       (\genblk2.pcpi_div_divisor [29]), .B
       (\genblk2.pcpi_div_dividend [29]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_49 ));
  NOR2BX1 \genblk2.pcpi_div_lte_2493_16_g1434 (.AN
       (\genblk2.pcpi_div_divisor [15]), .B
       (\genblk2.pcpi_div_dividend [15]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_48 ));
  NAND2BX1 \genblk2.pcpi_div_lte_2493_16_g1435 (.AN
       (\genblk2.pcpi_div_dividend [14]), .B
       (\genblk2.pcpi_div_divisor [14]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_47 ));
  NOR2BX1 \genblk2.pcpi_div_lte_2493_16_g1436 (.AN
       (\genblk2.pcpi_div_divisor [25]), .B
       (\genblk2.pcpi_div_dividend [25]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_46 ));
  NOR2BX1 \genblk2.pcpi_div_lte_2493_16_g1437 (.AN
       (\genblk2.pcpi_div_divisor [9]), .B
       (\genblk2.pcpi_div_dividend [9]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_44 ));
  NAND2BX1 \genblk2.pcpi_div_lte_2493_16_g1438 (.AN
       (\genblk2.pcpi_div_dividend [12]), .B
       (\genblk2.pcpi_div_divisor [12]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_43 ));
  NOR2BX1 \genblk2.pcpi_div_lte_2493_16_g1439 (.AN
       (\genblk2.pcpi_div_divisor [3]), .B
       (\genblk2.pcpi_div_dividend [3]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_42 ));
  NAND2BX1 \genblk2.pcpi_div_lte_2493_16_g1440 (.AN
       (\genblk2.pcpi_div_dividend [8]), .B
       (\genblk2.pcpi_div_divisor [8]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_41 ));
  NAND2BX1 \genblk2.pcpi_div_lte_2493_16_g1441 (.AN
       (\genblk2.pcpi_div_dividend [10]), .B
       (\genblk2.pcpi_div_divisor [10]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_40 ));
  NAND2BX1 \genblk2.pcpi_div_lte_2493_16_g1442 (.AN
       (\genblk2.pcpi_div_dividend [22]), .B
       (\genblk2.pcpi_div_divisor [22]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_39 ));
  NAND2BX1 \genblk2.pcpi_div_lte_2493_16_g1443 (.AN
       (\genblk2.pcpi_div_dividend [26]), .B
       (\genblk2.pcpi_div_divisor [26]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_38 ));
  NOR2BX1 \genblk2.pcpi_div_lte_2493_16_g1444 (.AN
       (\genblk2.pcpi_div_divisor [13]), .B
       (\genblk2.pcpi_div_dividend [13]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_37 ));
  NOR2BX1 \genblk2.pcpi_div_lte_2493_16_g1445 (.AN
       (\genblk2.pcpi_div_divisor [7]), .B
       (\genblk2.pcpi_div_dividend [7]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_36 ));
  NAND2BX1 \genblk2.pcpi_div_lte_2493_16_g1446 (.AN
       (\genblk2.pcpi_div_dividend [4]), .B
       (\genblk2.pcpi_div_divisor [4]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_35 ));
  NAND2BX1 \genblk2.pcpi_div_lte_2493_16_g1447 (.AN
       (\genblk2.pcpi_div_dividend [24]), .B
       (\genblk2.pcpi_div_divisor [24]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_34 ));
  NOR2BX1 \genblk2.pcpi_div_lte_2493_16_g1448 (.AN
       (\genblk2.pcpi_div_divisor [5]), .B
       (\genblk2.pcpi_div_dividend [5]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_33 ));
  NOR2BX1 \genblk2.pcpi_div_lte_2493_16_g1449 (.AN
       (\genblk2.pcpi_div_divisor [11]), .B
       (\genblk2.pcpi_div_dividend [11]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_32 ));
  NOR2BX1 \genblk2.pcpi_div_lte_2493_16_g1450 (.AN
       (\genblk2.pcpi_div_divisor [27]), .B
       (\genblk2.pcpi_div_dividend [27]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_31 ));
  NAND2BX1 \genblk2.pcpi_div_lte_2493_16_g1451 (.AN
       (\genblk2.pcpi_div_dividend [28]), .B
       (\genblk2.pcpi_div_divisor [28]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_30 ));
  NOR2BX1 \genblk2.pcpi_div_lte_2493_16_g1452 (.AN
       (\genblk2.pcpi_div_divisor [0]), .B
       (\genblk2.pcpi_div_dividend [0]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_45 ));
  INVX1 \genblk2.pcpi_div_lte_2493_16_g1453 (.A
       (\genblk2.pcpi_div_dividend [30]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_29 ));
  INVX1 \genblk2.pcpi_div_lte_2493_16_g1454 (.A
       (\genblk2.pcpi_div_dividend [7]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_28 ));
  INVX1 \genblk2.pcpi_div_lte_2493_16_g1455 (.A
       (\genblk2.pcpi_div_divisor [16]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_27 ));
  INVX1 \genblk2.pcpi_div_lte_2493_16_g1456 (.A
       (\genblk2.pcpi_div_divisor [6]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_26 ));
  INVX1 \genblk2.pcpi_div_lte_2493_16_g1457 (.A
       (\genblk2.pcpi_div_divisor [24]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_25 ));
  INVX1 \genblk2.pcpi_div_lte_2493_16_g1458 (.A
       (\genblk2.pcpi_div_dividend [17]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_24 ));
  INVX1 \genblk2.pcpi_div_lte_2493_16_g1459 (.A
       (\genblk2.pcpi_div_divisor [14]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_23 ));
  INVX1 \genblk2.pcpi_div_lte_2493_16_g1460 (.A
       (\genblk2.pcpi_div_divisor [2]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_22 ));
  INVX1 \genblk2.pcpi_div_lte_2493_16_g1461 (.A
       (\genblk2.pcpi_div_dividend [27]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_21 ));
  INVX1 \genblk2.pcpi_div_lte_2493_16_g1462 (.A
       (\genblk2.pcpi_div_dividend [21]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_20 ));
  INVX1 \genblk2.pcpi_div_lte_2493_16_g1463 (.A
       (\genblk2.pcpi_div_divisor [18]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_19 ));
  INVX1 \genblk2.pcpi_div_lte_2493_16_g1464 (.A
       (\genblk2.pcpi_div_divisor [8]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_18 ));
  INVX1 \genblk2.pcpi_div_lte_2493_16_g1465 (.A
       (\genblk2.pcpi_div_dividend [11]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_17 ));
  INVX1 \genblk2.pcpi_div_lte_2493_16_g1466 (.A
       (\genblk2.pcpi_div_divisor [12]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_16 ));
  INVX1 \genblk2.pcpi_div_lte_2493_16_g1467 (.A
       (\genblk2.pcpi_div_divisor [20]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_15 ));
  INVX1 \genblk2.pcpi_div_lte_2493_16_g1468 (.A
       (\genblk2.pcpi_div_dividend [3]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_14 ));
  INVX1 \genblk2.pcpi_div_lte_2493_16_g1469 (.A
       (\genblk2.pcpi_div_dividend [13]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_13 ));
  INVX1 \genblk2.pcpi_div_lte_2493_16_g1470 (.A
       (\genblk2.pcpi_div_divisor [26]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_12 ));
  INVX1 \genblk2.pcpi_div_lte_2493_16_g1471 (.A
       (\genblk2.pcpi_div_divisor [10]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_11 ));
  INVX1 \genblk2.pcpi_div_lte_2493_16_g1472 (.A
       (\genblk2.pcpi_div_divisor [4]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_10 ));
  INVX1 \genblk2.pcpi_div_lte_2493_16_g1473 (.A
       (\genblk2.pcpi_div_divisor [31]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_9 ));
  INVX1 \genblk2.pcpi_div_lte_2493_16_g1474 (.A
       (\genblk2.pcpi_div_divisor [22]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_8 ));
  INVX1 \genblk2.pcpi_div_lte_2493_16_g1475 (.A
       (\genblk2.pcpi_div_dividend [29]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_7 ));
  INVX1 \genblk2.pcpi_div_lte_2493_16_g1476 (.A
       (\genblk2.pcpi_div_dividend [9]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_6 ));
  INVX1 \genblk2.pcpi_div_lte_2493_16_g1477 (.A
       (\genblk2.pcpi_div_dividend [15]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_5 ));
  INVX1 \genblk2.pcpi_div_lte_2493_16_g1478 (.A
       (\genblk2.pcpi_div_divisor [28]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_4 ));
  INVX1 \genblk2.pcpi_div_lte_2493_16_g1479 (.A
       (\genblk2.pcpi_div_dividend [25]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_3 ));
  INVX1 \genblk2.pcpi_div_lte_2493_16_g1480 (.A
       (\genblk2.pcpi_div_dividend [19]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_2 ));
  INVX1 \genblk2.pcpi_div_lte_2493_16_g1481 (.A
       (\genblk2.pcpi_div_dividend [5]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_1 ));
  INVX1 \genblk2.pcpi_div_lte_2493_16_g1482 (.A
       (\genblk2.pcpi_div_dividend [23]), .Y
       (\genblk2.pcpi_div_lte_2493_16_n_0 ));
  CLKXOR2X1 g3(.A (n_6860), .B (inc_add_382_74_n_217), .Y (n_7126));
  CLKXOR2X1 g186397(.A (n_6853), .B (inc_add_382_74_n_252), .Y
       (n_7130));
  CLKXOR2X1 g186404(.A (n_6856), .B (inc_add_382_74_n_237), .Y
       (n_7137));
  CLKXOR2X1 g186406(.A (n_6850), .B (inc_add_382_74_n_267), .Y
       (n_7139));
  NAND2X1 g186411(.A (\reg_op2[0]_9669 ), .B (n_739), .Y (n_7145));
  MXI2XL g186412(.A (\reg_op1[31]_9668 ), .B (n_7146), .S0
       (\genblk2.pcpi_div_n_4742 ), .Y (n_7147));
  CLKXOR2X1 g186413(.A (\genblk2.pcpi_div_divisor [31]), .B
       (\genblk2.pcpi_div_dividend [31]), .Y (n_7146));
  BUFX20 fopt186769(.A (\reg_op2[27]_9696 ), .Y (pcpi_rs2[27]));
  BUFX20 fopt186774(.A (\reg_op2[23]_9692 ), .Y (pcpi_rs2[23]));
  BUFX20 fopt186779(.A (\reg_op2[25]_9694 ), .Y (pcpi_rs2[25]));
  BUFX20 fopt186784(.A (\reg_op2[29]_9698 ), .Y (pcpi_rs2[29]));
  BUFX20 fopt186789(.A (\reg_op1[4]_9641 ), .Y (pcpi_rs1[4]));
  BUFX20 fopt186794(.A (\reg_op2[30]_9699 ), .Y (pcpi_rs2[30]));
  BUFX20 fopt186799(.A (\reg_op1[27]_9664 ), .Y (pcpi_rs1[27]));
  BUFX20 fopt186804(.A (\reg_op1[20]_9657 ), .Y (pcpi_rs1[20]));
  BUFX20 fopt186809(.A (\reg_op1[21]_9658 ), .Y (pcpi_rs1[21]));
  BUFX20 fopt186814(.A (\reg_op1[22]_9659 ), .Y (pcpi_rs1[22]));
  BUFX20 fopt186819(.A (\reg_op1[23]_9660 ), .Y (pcpi_rs1[23]));
  BUFX20 fopt186824(.A (\reg_op1[24]_9661 ), .Y (pcpi_rs1[24]));
  BUFX20 fopt186829(.A (\reg_op2[3]_9672 ), .Y (mem_la_wdata[3]));
  BUFX20 fopt186834(.A (\reg_op1[25]_9662 ), .Y (pcpi_rs1[25]));
  BUFX20 fopt186839(.A (\reg_op1[26]_9663 ), .Y (pcpi_rs1[26]));
  BUFX20 fopt186844(.A (\reg_op1[28]_9665 ), .Y (pcpi_rs1[28]));
  BUFX20 fopt186849(.A (\reg_op2[20]_9689 ), .Y (pcpi_rs2[20]));
  BUFX20 fopt186854(.A (\reg_op1[29]_9666 ), .Y (pcpi_rs1[29]));
  BUFX20 fopt186859(.A (\reg_op1[30]_9667 ), .Y (pcpi_rs1[30]));
  BUFX20 fopt186864(.A (\reg_op1[17]_9654 ), .Y (pcpi_rs1[17]));
  BUFX20 fopt186869(.A (\reg_op2[4]_9673 ), .Y (pcpi_rs2[4]));
  BUFX20 fopt186874(.A (\reg_op1[18]_9655 ), .Y (pcpi_rs1[18]));
  BUFX20 fopt186879(.A (\reg_op1[19]_9656 ), .Y (pcpi_rs1[19]));
  BUFX20 fopt186884(.A (\reg_op2[24]_9693 ), .Y (pcpi_rs2[24]));
  BUFX20 fopt186889(.A (\reg_op2[26]_9695 ), .Y (pcpi_rs2[26]));
  BUFX20 fopt186894(.A (\reg_op2[28]_9697 ), .Y (pcpi_rs2[28]));
  BUFX20 fopt186899(.A (\reg_op1[31]_9668 ), .Y (pcpi_rs1[31]));
  BUFX20 fopt186904(.A (\reg_op2[22]_9691 ), .Y (pcpi_rs2[22]));
  BUFX20 fopt186909(.A (\reg_op2[3]_9672 ), .Y (pcpi_rs2[3]));
  BUFX20 fopt186914(.A (\reg_op2[31]_9700 ), .Y (pcpi_rs2[31]));
  BUFX20 fopt186929(.A (\reg_op2[6]_9675 ), .Y (mem_la_wdata[6]));
  BUFX20 fopt186934(.A (\reg_op1[9]_9646 ), .Y (pcpi_rs1[9]));
  BUFX20 fopt186939(.A (\reg_op1[11]_9648 ), .Y (pcpi_rs1[11]));
  BUFX20 fopt186944(.A (\reg_op1[12]_9649 ), .Y (pcpi_rs1[12]));
  BUFX20 fopt186949(.A (\reg_op2[15]_9684 ), .Y (pcpi_rs2[15]));
  BUFX20 fopt186954(.A (\reg_op1[10]_9647 ), .Y (pcpi_rs1[10]));
  BUFX20 fopt186959(.A (\reg_op2[9]_9678 ), .Y (pcpi_rs2[9]));
  BUFX20 fopt186964(.A (\reg_op2[10]_9679 ), .Y (pcpi_rs2[10]));
  BUFX20 fopt186969(.A (\reg_op2[16]_9685 ), .Y (pcpi_rs2[16]));
  BUFX20 fopt186974(.A (\reg_op2[14]_9683 ), .Y (pcpi_rs2[14]));
  BUFX20 fopt186979(.A (\reg_op2[19]_9688 ), .Y (pcpi_rs2[19]));
  BUFX20 fopt186984(.A (\reg_op2[11]_9680 ), .Y (pcpi_rs2[11]));
  BUFX20 fopt186989(.A (\reg_op2[12]_9681 ), .Y (pcpi_rs2[12]));
  BUFX20 fopt186994(.A (\reg_op2[13]_9682 ), .Y (pcpi_rs2[13]));
  BUFX20 fopt186999(.A (\reg_op2[18]_9687 ), .Y (pcpi_rs2[18]));
  BUFX20 fopt187004(.A (\reg_op2[17]_9686 ), .Y (pcpi_rs2[17]));
  BUFX20 fopt187009(.A (\reg_op2[2]_9671 ), .Y (pcpi_rs2[2]));
  BUFX20 fopt187014(.A (\reg_op2[7]_9676 ), .Y (mem_la_wdata[7]));
  BUFX20 fopt187019(.A (\reg_op2[4]_9673 ), .Y (mem_la_wdata[4]));
  BUFX20 fopt187024(.A (\reg_op1[15]_9652 ), .Y (pcpi_rs1[15]));
  BUFX20 fopt187029(.A (\reg_op2[6]_9675 ), .Y (pcpi_rs2[6]));
  BUFX20 fopt187034(.A (\reg_op1[2]_9639 ), .Y (pcpi_rs1[2]));
  BUFX20 fopt187039(.A (\reg_op1[13]_9650 ), .Y (pcpi_rs1[13]));
  BUFX20 fopt187044(.A (\reg_op2[8]_9677 ), .Y (pcpi_rs2[8]));
  BUFX20 fopt187049(.A (\reg_op2[1]_9670 ), .Y (mem_la_wdata[1]));
  BUFX20 fopt187054(.A (mem_valid_9465), .Y (mem_valid));
  BUFX20 fopt187059(.A (\reg_op2[5]_9674 ), .Y (pcpi_rs2[5]));
  BUFX20 fopt187064(.A (\reg_op2[21]_9690 ), .Y (pcpi_rs2[21]));
  BUFX20 fopt187069(.A (\reg_op2[1]_9670 ), .Y (pcpi_rs2[1]));
  BUFX20 fopt187074(.A (reg_op1[0]), .Y (pcpi_rs1[0]));
  BUFX20 fopt187079(.A (\reg_op1[16]_9653 ), .Y (pcpi_rs1[16]));
  BUFX20 fopt187084(.A (\reg_op2[0]_9669 ), .Y (pcpi_rs2[0]));
  BUFX20 fopt187089(.A (\reg_op1[14]_9651 ), .Y (pcpi_rs1[14]));
  BUFX20 fopt187094(.A (\reg_op2[2]_9671 ), .Y (mem_la_wdata[2]));
  BUFX20 fopt187099(.A (\reg_op1[7]_9644 ), .Y (pcpi_rs1[7]));
  BUFX20 fopt187104(.A (\reg_op1[5]_9642 ), .Y (pcpi_rs1[5]));
  BUFX20 fopt187109(.A (\reg_op2[7]_9676 ), .Y (pcpi_rs2[7]));
  BUFX20 fopt187114(.A (\reg_op1[3]_9640 ), .Y (pcpi_rs1[3]));
  BUFX20 fopt187119(.A (\reg_op2[5]_9674 ), .Y (mem_la_wdata[5]));
  BUFX20 fopt187124(.A (\reg_op1[1]_9638 ), .Y (pcpi_rs1[1]));
  BUFX20 fopt187129(.A (\reg_op1[8]_9645 ), .Y (pcpi_rs1[8]));
  BUFX20 fopt187134(.A (\reg_op1[6]_9643 ), .Y (pcpi_rs1[6]));
  BUFX20 fopt187139(.A (\reg_op2[0]_9669 ), .Y (mem_la_wdata[0]));
  NOR3BXL g82728__187171(.AN (n_5599), .B (n_6530), .C (n_5598), .Y
       (n_8138));
  NOR4BBX1 g82731__187322(.AN (n_5610), .BN (n_5590), .C (n_5611), .D
       (n_5591), .Y (n_8325));
  BUFX20 fopt187452(.A (n_8490), .Y (mem_la_addr[29]));
  MXI2XL g187453(.A (n_716), .B (n_7126), .S0 (n_313), .Y (n_8490));
  MX2X1 g187454(.A (n_8490), .B (n_5689), .S0 (n_472), .Y (n_8493));
  BUFX20 fopt187468(.A (n_11855), .Y (mem_la_addr[28]));
  MX2X1 g187470(.A (n_11855), .B (n_5688), .S0 (n_472), .Y (n_8514));
  BUFX20 fopt187484(.A (n_11833), .Y (mem_la_addr[27]));
  MX2X1 g187486(.A (n_11833), .B (n_5687), .S0 (n_472), .Y (n_8535));
  BUFX20 fopt187500(.A (n_8553), .Y (mem_la_addr[18]));
  MX2XL g187501(.A (\reg_op1[18]_9655 ), .B (n_6819), .S0 (n_313), .Y
       (n_8553));
  MX2X1 g187502(.A (n_8553), .B (n_5678), .S0 (n_472), .Y (n_8556));
  BUFX20 fopt187516(.A (n_11834), .Y (mem_la_addr[26]));
  MX2X1 g187518(.A (n_11834), .B (n_5686), .S0 (n_472), .Y (n_8577));
  BUFX20 fopt187532(.A (n_8595), .Y (mem_la_addr[25]));
  MXI2XL g187533(.A (n_5784), .B (n_7137), .S0 (n_313), .Y (n_8595));
  MX2X1 g187534(.A (n_8595), .B (n_5685), .S0 (n_472), .Y (n_8598));
  BUFX20 fopt187548(.A (n_11857), .Y (mem_la_addr[24]));
  MX2X1 g187550(.A (n_11857), .B (n_5684), .S0 (n_472), .Y (n_8619));
  BUFX20 fopt187564(.A (n_11836), .Y (mem_la_addr[23]));
  MX2X1 g187566(.A (n_11836), .B (n_5683), .S0 (n_472), .Y (n_8640));
  BUFX20 fopt187580(.A (n_8658), .Y (mem_la_addr[22]));
  MXI2XL g187581(.A (n_576), .B (n_7130), .S0 (n_313), .Y (n_8658));
  MX2X1 g187582(.A (n_8658), .B (n_5682), .S0 (n_472), .Y (n_8661));
  BUFX20 fopt187596(.A (n_11859), .Y (mem_la_addr[21]));
  MX2X1 g187598(.A (n_11859), .B (n_5681), .S0 (n_472), .Y (n_8682));
  BUFX20 fopt187612(.A (n_11838), .Y (mem_la_addr[20]));
  MX2X1 g187614(.A (n_11838), .B (n_5680), .S0 (n_472), .Y (n_8703));
  BUFX20 fopt187628(.A (n_8721), .Y (mem_la_addr[19]));
  MXI2XL g187629(.A (n_747), .B (n_7139), .S0 (n_313), .Y (n_8721));
  MX2X1 g187630(.A (n_8721), .B (n_5679), .S0 (n_472), .Y (n_8724));
  BUFX20 fopt187644(.A (n_11861), .Y (mem_la_addr[17]));
  MX2X1 g187646(.A (n_11861), .B (n_5677), .S0 (n_472), .Y (n_8745));
  BUFX20 fopt187660(.A (n_11840), .Y (mem_la_addr[16]));
  MX2X1 g187662(.A (n_11840), .B (n_5676), .S0 (n_472), .Y (n_8766));
  BUFX20 fopt187676(.A (n_8784), .Y (mem_la_addr[15]));
  MX2XL g187677(.A (\reg_op1[15]_9652 ), .B (n_6816), .S0 (n_313), .Y
       (n_8784));
  MX2X1 g187678(.A (n_8784), .B (n_5675), .S0 (n_472), .Y (n_8787));
  BUFX20 fopt187692(.A (n_11863), .Y (mem_la_addr[30]));
  MX2X1 g187694(.A (n_11863), .B (n_5690), .S0 (n_472), .Y (n_8808));
  BUFX20 fopt187708(.A (n_11842), .Y (mem_la_addr[2]));
  MX2X1 g187710(.A (n_11842), .B (n_5662), .S0 (n_472), .Y (n_8829));
  BUFX20 fopt187724(.A (n_8847), .Y (mem_la_addr[13]));
  MX2XL g187725(.A (\reg_op1[13]_9650 ), .B (n_6814), .S0 (n_313), .Y
       (n_8847));
  MX2X1 g187726(.A (n_8847), .B (n_5673), .S0 (n_472), .Y (n_8850));
  BUFX20 fopt187740(.A (n_8868), .Y (mem_la_addr[12]));
  MX2XL g187741(.A (\reg_op1[12]_9649 ), .B (n_6813), .S0 (n_313), .Y
       (n_8868));
  MX2X1 g187742(.A (n_8868), .B (n_5672), .S0 (n_472), .Y (n_8871));
  BUFX20 fopt187756(.A (n_11843), .Y (mem_la_wdata[10]));
  MX2X1 g187758(.A (n_11843), .B (n_5640), .S0 (n_542), .Y (n_8892));
  BUFX20 fopt187772(.A (n_8910), .Y (mem_la_addr[11]));
  MX2XL g187773(.A (\reg_op1[11]_9648 ), .B (n_6812), .S0 (n_313), .Y
       (n_8910));
  MX2X1 g187774(.A (n_8910), .B (n_5671), .S0 (n_472), .Y (n_8913));
  BUFX20 fopt187788(.A (n_8931), .Y (mem_la_addr[9]));
  MX2XL g187789(.A (\reg_op1[9]_9646 ), .B (n_6810), .S0 (n_313), .Y
       (n_8931));
  MX2X1 g187790(.A (n_8931), .B (n_5669), .S0 (n_472), .Y (n_8934));
  BUFX20 fopt187804(.A (n_8952), .Y (mem_la_addr[8]));
  MX2XL g187805(.A (\reg_op1[8]_9645 ), .B (n_6809), .S0 (n_313), .Y
       (n_8952));
  MX2X1 g187806(.A (n_8952), .B (n_5668), .S0 (n_472), .Y (n_8955));
  BUFX20 fopt187820(.A (n_11844), .Y (mem_la_wdata[14]));
  MX2X1 g187822(.A (n_11844), .B (n_5644), .S0 (n_542), .Y (n_8976));
  BUFX20 fopt187836(.A (n_8994), .Y (mem_la_addr[7]));
  MX2XL g187837(.A (\reg_op1[7]_9644 ), .B (n_6808), .S0 (n_313), .Y
       (n_8994));
  MX2X1 g187838(.A (n_8994), .B (n_5667), .S0 (n_472), .Y (n_8997));
  BUFX20 fopt187852(.A (n_11845), .Y (mem_la_addr[5]));
  MX2X1 g187854(.A (n_11845), .B (n_5665), .S0 (n_472), .Y (n_9018));
  BUFX20 fopt187868(.A (n_11846), .Y (mem_la_addr[4]));
  MX2X1 g187870(.A (n_11846), .B (n_5664), .S0 (n_472), .Y (n_9039));
  BUFX20 fopt187884(.A (n_11847), .Y (mem_la_addr[3]));
  MX2X1 g187886(.A (n_11847), .B (n_5663), .S0 (n_472), .Y (n_9060));
  BUFX20 fopt187900(.A (n_9078), .Y (mem_la_wstrb[3]));
  OR2X1 g89840__187901(.A (n_608), .B (n_6222), .Y (n_9078));
  AO22X1 g187902(.A0 (n_9078), .A1 (n_2150), .B0 (n_5629), .B1
       (n_1950), .Y (n_9081));
  BUFX20 fopt187916(.A (n_9099), .Y (mem_la_wstrb[2]));
  OR2X1 g89825__187917(.A (n_608), .B (n_340), .Y (n_9099));
  AO22X1 g187918(.A0 (n_9099), .A1 (n_2150), .B0 (n_5628), .B1
       (n_1950), .Y (n_9102));
  BUFX20 fopt187932(.A (n_9120), .Y (mem_la_wstrb[1]));
  OR2X1 g89900__187933(.A (n_6082), .B (n_657), .Y (n_9120));
  AO22X1 g187934(.A0 (n_9120), .A1 (n_2150), .B0 (n_5627), .B1
       (n_1950), .Y (n_9123));
  BUFX20 fopt187948(.A (n_9141), .Y (mem_la_wstrb[0]));
  OR2X1 g89906__187949(.A (n_6082), .B (n_6122), .Y (n_9141));
  AO22X1 g187950(.A0 (n_9141), .A1 (n_2150), .B0 (n_5626), .B1
       (n_1950), .Y (n_9144));
  BUFX20 fopt187964(.A (n_9162), .Y (mem_la_wdata[16]));
  OR2X1 g90004__187965(.A (n_6115), .B (n_6113), .Y (n_9162));
  MX2X1 g187966(.A (n_9162), .B (n_5646), .S0 (n_542), .Y (n_9165));
  BUFX20 fopt187980(.A (n_9183), .Y (mem_la_wdata[23]));
  OR2X1 g89998__187981(.A (n_6119), .B (n_6118), .Y (n_9183));
  MX2X1 g187982(.A (n_9183), .B (n_5653), .S0 (n_542), .Y (n_9186));
  BUFX20 fopt187996(.A (n_9204), .Y (mem_la_wdata[20]));
  OR2X1 g90001__187997(.A (n_6072), .B (n_6110), .Y (n_9204));
  MX2X1 g187998(.A (n_9204), .B (n_5650), .S0 (n_542), .Y (n_9207));
  BUFX20 fopt188012(.A (n_9225), .Y (mem_la_wdata[18]));
  OR2X1 g90003__188013(.A (n_6070), .B (n_6121), .Y (n_9225));
  MX2X1 g188014(.A (n_9225), .B (n_5648), .S0 (n_542), .Y (n_9228));
  BUFX20 fopt188028(.A (n_9246), .Y (mem_la_wdata[22]));
  OR2X1 g89999__188029(.A (n_6114), .B (n_6112), .Y (n_9246));
  MX2X1 g188030(.A (n_9246), .B (n_5652), .S0 (n_542), .Y (n_9249));
  BUFX20 fopt188044(.A (n_9267), .Y (mem_la_wdata[29]));
  OR2X1 g89833__188045(.A (n_6098), .B (n_11765), .Y (n_9267));
  MX2X1 g188046(.A (n_9267), .B (n_5659), .S0 (n_542), .Y (n_9270));
  BUFX20 fopt188060(.A (n_9288), .Y (mem_la_wdata[24]));
  OR2X1 g89842__188061(.A (n_6134), .B (n_11759), .Y (n_9288));
  MX2X1 g188062(.A (n_9288), .B (n_5654), .S0 (n_542), .Y (n_9291));
  BUFX20 fopt188076(.A (n_9309), .Y (mem_la_wdata[27]));
  OR2X1 g89834__188077(.A (n_6101), .B (n_11762), .Y (n_9309));
  MX2X1 g188078(.A (n_9309), .B (n_5657), .S0 (n_542), .Y (n_9312));
  BUFX20 fopt188092(.A (n_9330), .Y (mem_la_wdata[26]));
  OR2X1 g89835__188093(.A (n_6103), .B (n_11764), .Y (n_9330));
  MX2X1 g188094(.A (n_9330), .B (n_5656), .S0 (n_542), .Y (n_9333));
  BUFX20 fopt188108(.A (n_9351), .Y (mem_la_addr[6]));
  MX2XL g188109(.A (\reg_op1[6]_9643 ), .B (n_6807), .S0 (n_313), .Y
       (n_9351));
  MX2X1 g188110(.A (n_9351), .B (n_5666), .S0 (n_472), .Y (n_9354));
  BUFX20 fopt188124(.A (n_9372), .Y (mem_la_wdata[30]));
  OR2X1 g89823__188125(.A (n_6141), .B (n_11761), .Y (n_9372));
  MX2X1 g188126(.A (n_9372), .B (n_5660), .S0 (n_542), .Y (n_9375));
  BUFX20 fopt188140(.A (n_9393), .Y (mem_la_wdata[31]));
  OR2X1 g89838__188141(.A (n_6105), .B (n_11763), .Y (n_9393));
  MX2X1 g188142(.A (n_9393), .B (n_5661), .S0 (n_542), .Y (n_9396));
  BUFX20 fopt188156(.A (n_9414), .Y (mem_la_addr[14]));
  MX2XL g188157(.A (\reg_op1[14]_9651 ), .B (n_6815), .S0 (n_313), .Y
       (n_9414));
  MX2X1 g188158(.A (n_9414), .B (n_5674), .S0 (n_472), .Y (n_9417));
  BUFX20 fopt188172(.A (n_9435), .Y (mem_la_addr[10]));
  MX2XL g188173(.A (\reg_op1[10]_9647 ), .B (n_6811), .S0 (n_313), .Y
       (n_9435));
  MX2X1 g188174(.A (n_9435), .B (n_5670), .S0 (n_472), .Y (n_9438));
  BUFX20 fopt188188(.A (n_9456), .Y (mem_la_wdata[28]));
  OR2X1 g89841__188189(.A (n_6104), .B (n_11760), .Y (n_9456));
  MX2X1 g188190(.A (n_9456), .B (n_5658), .S0 (n_542), .Y (n_9459));
  BUFX20 fopt188204(.A (n_9477), .Y (mem_la_wdata[25]));
  OR2X1 g89837__188205(.A (n_6097), .B (n_11766), .Y (n_9477));
  MX2X1 g188206(.A (n_9477), .B (n_5655), .S0 (n_542), .Y (n_9480));
  BUFX20 fopt188220(.A (n_9498), .Y (mem_la_wdata[19]));
  OR2X1 g90002__188221(.A (n_6071), .B (n_6117), .Y (n_9498));
  MX2X1 g188222(.A (n_9498), .B (n_5649), .S0 (n_542), .Y (n_9501));
  BUFX20 fopt188236(.A (n_9519), .Y (mem_la_wdata[21]));
  OR2X1 g90000__188237(.A (n_6073), .B (n_6106), .Y (n_9519));
  MX2X1 g188238(.A (n_9519), .B (n_5651), .S0 (n_542), .Y (n_9522));
  BUFX20 fopt188252(.A (n_9540), .Y (mem_la_wdata[17]));
  OR2X1 g89955__188253(.A (n_6124), .B (n_6111), .Y (n_9540));
  MX2X1 g188254(.A (n_9540), .B (n_5647), .S0 (n_542), .Y (n_9543));
  BUFX20 fopt188268(.A (n_11848), .Y (mem_la_wdata[15]));
  MX2X1 g188270(.A (n_11848), .B (n_5645), .S0 (n_542), .Y (n_9564));
  BUFX20 fopt188284(.A (n_11849), .Y (mem_la_wdata[13]));
  MX2X1 g188286(.A (n_11849), .B (n_5643), .S0 (n_542), .Y (n_9585));
  BUFX20 fopt188300(.A (n_11850), .Y (mem_la_wdata[12]));
  MX2X1 g188302(.A (n_11850), .B (n_5642), .S0 (n_542), .Y (n_9606));
  BUFX20 fopt188316(.A (n_11851), .Y (mem_la_wdata[11]));
  MX2X1 g188318(.A (n_11851), .B (n_5641), .S0 (n_542), .Y (n_9627));
  BUFX20 fopt188332(.A (n_11852), .Y (mem_la_wdata[9]));
  MX2X1 g188334(.A (n_11852), .B (n_5639), .S0 (n_542), .Y (n_9648));
  BUFX20 fopt188348(.A (n_11853), .Y (mem_la_wdata[8]));
  MX2X1 g188350(.A (n_11853), .B (n_5638), .S0 (n_542), .Y (n_9669));
  BUFX20 fopt188364(.A (n_9687), .Y (mem_la_addr[31]));
  MX2XL g188365(.A (\reg_op1[31]_9668 ), .B (n_6832), .S0 (n_313), .Y
       (n_9687));
  MX2X1 g188366(.A (n_9687), .B (n_5691), .S0 (n_472), .Y (n_9690));
  BUFX20 drc188629(.A (n_5597), .Y (pcpi_insn[12]));
  BUFX20 drc188644(.A (n_5599), .Y (pcpi_insn[14]));
  BUFX20 drc188659(.A (n_5598), .Y (pcpi_insn[13]));
  BUFX20 fopt188674(.A (n_5587), .Y (pcpi_insn[2]));
  BUFX20 fopt188689(.A (n_5588), .Y (pcpi_insn[3]));
  BUFX20 fopt188704(.A (n_5589), .Y (pcpi_insn[4]));
  BUFX20 fopt188719(.A (n_5590), .Y (pcpi_insn[5]));
  BUFX20 fopt188734(.A (n_5591), .Y (pcpi_insn[6]));
  BUFX20 fopt188749(.A (n_5586), .Y (pcpi_insn[1]));
  NOR4BBX1 g82732__188750(.AN (n_5589), .BN (n_5586), .C (n_5588), .D
       (n_5587), .Y (n_10451));
  BUFX20 fopt188764(.A (n_5585), .Y (pcpi_insn[0]));
  BUFX20 fopt188779(.A (n_5610), .Y (pcpi_insn[25]));
  NAND4BXL g90105__188780(.AN (n_5591), .B (n_5589), .C (n_5590), .D
       (n_5610), .Y (n_10491));
  BUFX20 fopt188794(.A (n_5611), .Y (pcpi_insn[26]));
  BUFX20 fopt188809(.A (n_5612), .Y (pcpi_insn[27]));
  NOR4X1 g90109__188810(.A (n_5612), .B (n_5611), .C (n_5613), .D
       (n_5614), .Y (n_10531));
  BUFX20 fopt188824(.A (n_5613), .Y (pcpi_insn[28]));
  NOR4X1 g82733__188825(.A (n_5613), .B (n_5612), .C (n_5614), .D
       (n_5615), .Y (n_10551));
  BUFX20 fopt188839(.A (n_5616), .Y (pcpi_insn[31]));
  BUFX20 fopt188854(.A (n_5614), .Y (pcpi_insn[29]));
  BUFX20 fopt188869(.A (n_5615), .Y (pcpi_insn[30]));
  BUFX20 fopt188884(.A (n_5617), .Y (pcpi_valid));
  EDFFX2 \genblk2.pcpi_div_outsign_reg (.CK (clk), .D (n_5262), .E
       (n_668), .Q (\genblk2.pcpi_div_outsign ), .QN (n_5994));
  DFFX2 instr_rdinstrh_reg(.CK (clk), .D (n_5103), .Q (instr_rdinstrh),
       .QN (n_558));
  DFFX2 \cpu_state_reg[5] (.CK (clk), .D (n_5037), .Q (cpu_state[5]),
       .QN (n_548));
  DFFX2 instr_sub_reg(.CK (clk), .D (n_2950), .Q (instr_sub), .QN
       (sub_1235_38_Y_add_1235_58_n_1443));
  DFFX2 \genblk1.pcpi_mul_rs2_reg[32] (.CK (clk), .D (n_2010), .Q
       (\genblk1.pcpi_mul_rs2 [32]), .QN
       (\genblk1.pcpi_mul_mul_2366_47_n_172 ));
  DFFX1 \genblk1.pcpi_mul_rs1_reg[24] (.CK (clk), .D (n_1695), .Q
       (\genblk1.pcpi_mul_rs1 [24]), .QN
       (\genblk1.pcpi_mul_mul_2366_47_n_99 ));
  DFFX1 \genblk1.pcpi_mul_rs1_reg[15] (.CK (clk), .D (n_1701), .Q
       (\genblk1.pcpi_mul_rs1 [15]), .QN
       (\genblk1.pcpi_mul_mul_2366_47_n_97 ));
  DFFX1 \genblk1.pcpi_mul_rs1_reg[22] (.CK (clk), .D (n_1696), .Q
       (\genblk1.pcpi_mul_rs1 [22]), .QN
       (\genblk1.pcpi_mul_mul_2366_47_n_95 ));
  DFFX1 \genblk1.pcpi_mul_rs1_reg[3] (.CK (clk), .D (n_1707), .Q
       (\genblk1.pcpi_mul_rs1 [3]), .QN
       (\genblk1.pcpi_mul_mul_2366_47_n_93 ));
  DFFX1 \genblk1.pcpi_mul_rs1_reg[7] (.CK (clk), .D (n_1672), .Q
       (\genblk1.pcpi_mul_rs1 [7]), .QN
       (\genblk1.pcpi_mul_mul_2366_47_n_91 ));
  DFFX1 \genblk1.pcpi_mul_rs1_reg[16] (.CK (clk), .D (n_1668), .Q
       (\genblk1.pcpi_mul_rs1 [16]), .QN
       (\genblk1.pcpi_mul_mul_2366_47_n_89 ));
  DFFX1 \genblk1.pcpi_mul_rs1_reg[20] (.CK (clk), .D (n_1667), .Q
       (\genblk1.pcpi_mul_rs1 [20]), .QN
       (\genblk1.pcpi_mul_mul_2366_47_n_87 ));
  DFFX1 \genblk1.pcpi_mul_rs1_reg[8] (.CK (clk), .D (n_1705), .Q
       (\genblk1.pcpi_mul_rs1 [8]), .QN
       (\genblk1.pcpi_mul_mul_2366_47_n_85 ));
  DFFX1 \genblk1.pcpi_mul_rs1_reg[17] (.CK (clk), .D (n_1662), .Q
       (\genblk1.pcpi_mul_rs1 [17]), .QN
       (\genblk1.pcpi_mul_mul_2366_47_n_83 ));
  DFFX1 \genblk1.pcpi_mul_rs1_reg[1] (.CK (clk), .D (n_1691), .Q
       (\genblk1.pcpi_mul_rs1 [1]), .QN
       (\genblk1.pcpi_mul_mul_2366_47_n_81 ));
  DFFX1 \genblk1.pcpi_mul_rs1_reg[18] (.CK (clk), .D (n_1699), .Q
       (\genblk1.pcpi_mul_rs1 [18]), .QN
       (\genblk1.pcpi_mul_mul_2366_47_n_79 ));
  DFFX1 \genblk1.pcpi_mul_rs1_reg[27] (.CK (clk), .D (n_1693), .Q
       (\genblk1.pcpi_mul_rs1 [27]), .QN
       (\genblk1.pcpi_mul_mul_2366_47_n_77 ));
  DFFX1 \genblk1.pcpi_mul_rs1_reg[9] (.CK (clk), .D (n_1704), .Q
       (\genblk1.pcpi_mul_rs1 [9]), .QN
       (\genblk1.pcpi_mul_mul_2366_47_n_75 ));
  DFFX1 \genblk1.pcpi_mul_rs1_reg[19] (.CK (clk), .D (n_1698), .Q
       (\genblk1.pcpi_mul_rs1 [19]), .QN
       (\genblk1.pcpi_mul_mul_2366_47_n_73 ));
  DFFX1 \genblk1.pcpi_mul_rs1_reg[4] (.CK (clk), .D (n_1669), .Q
       (\genblk1.pcpi_mul_rs1 [4]), .QN
       (\genblk1.pcpi_mul_mul_2366_47_n_71 ));
  DFFX1 \genblk1.pcpi_mul_rs1_reg[10] (.CK (clk), .D (n_1700), .Q
       (\genblk1.pcpi_mul_rs1 [10]), .QN
       (\genblk1.pcpi_mul_mul_2366_47_n_69 ));
  DFFX1 \genblk1.pcpi_mul_rs1_reg[21] (.CK (clk), .D (n_1697), .Q
       (\genblk1.pcpi_mul_rs1 [21]), .QN
       (\genblk1.pcpi_mul_mul_2366_47_n_67 ));
  DFFX1 \genblk1.pcpi_mul_rs1_reg[28] (.CK (clk), .D (n_1666), .Q
       (\genblk1.pcpi_mul_rs1 [28]), .QN
       (\genblk1.pcpi_mul_mul_2366_47_n_65 ));
  DFFX1 \genblk1.pcpi_mul_rs1_reg[30] (.CK (clk), .D (n_1692), .Q
       (\genblk1.pcpi_mul_rs1 [30]), .QN
       (\genblk1.pcpi_mul_mul_2366_47_n_63 ));
  DFFX1 \genblk1.pcpi_mul_rs1_reg[29] (.CK (clk), .D (n_1665), .Q
       (\genblk1.pcpi_mul_rs1 [29]), .QN
       (\genblk1.pcpi_mul_mul_2366_47_n_61 ));
  DFFX1 \genblk1.pcpi_mul_rs1_reg[6] (.CK (clk), .D (n_1677), .Q
       (\genblk1.pcpi_mul_rs1 [6]), .QN
       (\genblk1.pcpi_mul_mul_2366_47_n_59 ));
  DFFX1 \genblk1.pcpi_mul_rs1_reg[2] (.CK (clk), .D (n_1708), .Q
       (\genblk1.pcpi_mul_rs1 [2]), .QN
       (\genblk1.pcpi_mul_mul_2366_47_n_57 ));
  DFFX1 \genblk1.pcpi_mul_rs1_reg[26] (.CK (clk), .D (n_1675), .Q
       (\genblk1.pcpi_mul_rs1 [26]), .QN
       (\genblk1.pcpi_mul_mul_2366_47_n_55 ));
  DFFX1 \genblk1.pcpi_mul_rs1_reg[25] (.CK (clk), .D (n_1694), .Q
       (\genblk1.pcpi_mul_rs1 [25]), .QN
       (\genblk1.pcpi_mul_mul_2366_47_n_53 ));
  DFFX1 \genblk1.pcpi_mul_rs1_reg[11] (.CK (clk), .D (n_1670), .Q
       (\genblk1.pcpi_mul_rs1 [11]), .QN
       (\genblk1.pcpi_mul_mul_2366_47_n_51 ));
  DFFX1 \genblk1.pcpi_mul_rs1_reg[23] (.CK (clk), .D (n_1678), .Q
       (\genblk1.pcpi_mul_rs1 [23]), .QN
       (\genblk1.pcpi_mul_mul_2366_47_n_49 ));
  DFFX1 \genblk1.pcpi_mul_rs1_reg[5] (.CK (clk), .D (n_1706), .Q
       (\genblk1.pcpi_mul_rs1 [5]), .QN
       (\genblk1.pcpi_mul_mul_2366_47_n_47 ));
  DFFX1 \genblk1.pcpi_mul_rs1_reg[12] (.CK (clk), .D (n_1703), .Q
       (\genblk1.pcpi_mul_rs1 [12]), .QN
       (\genblk1.pcpi_mul_mul_2366_47_n_45 ));
  DFFX1 \genblk1.pcpi_mul_rs1_reg[31] (.CK (clk), .D (n_1663), .Q
       (\genblk1.pcpi_mul_rs1 [31]), .QN
       (\genblk1.pcpi_mul_mul_2366_47_n_43 ));
  DFFX1 \genblk1.pcpi_mul_rs1_reg[13] (.CK (clk), .D (n_1676), .Q
       (\genblk1.pcpi_mul_rs1 [13]), .QN
       (\genblk1.pcpi_mul_mul_2366_47_n_41 ));
  DFFX1 \genblk1.pcpi_mul_rs1_reg[14] (.CK (clk), .D (n_1702), .Q
       (\genblk1.pcpi_mul_rs1 [14]), .QN
       (\genblk1.pcpi_mul_mul_2366_47_n_39 ));
  DFFX1 \genblk1.pcpi_mul_rs1_reg[32] (.CK (clk), .D (n_2262), .Q
       (\genblk1.pcpi_mul_rs1 [32]), .QN
       (\genblk1.pcpi_mul_mul_2366_47_n_37 ));
  DFFX1 \genblk1.pcpi_mul_rs2_reg[0] (.CK (clk), .D (n_1679), .Q
       (\genblk1.pcpi_mul_rs2 [0]), .QN
       (\genblk1.pcpi_mul_mul_2366_47_n_35 ));
  NOR2BX4 g2(.AN (pcpi_ready), .B (n_356), .Y (n_11689));
  NOR2BX4 g189415(.AN (\genblk1.pcpi_mul_shift_out ), .B (n_6527), .Y
       (n_11690));
  NOR2BX1 g189416(.AN (n_6059), .B (n_6051), .Y (n_11691));
  MXI2XL g189417(.A (\genblk2.pcpi_div_dividend [14]), .B
       (\genblk2.pcpi_div_quotient [14]), .S0 (\genblk2.pcpi_div_n_2109
       ), .Y (n_11692));
  MXI2XL g189418(.A (\genblk2.pcpi_div_dividend [10]), .B
       (\genblk2.pcpi_div_quotient [10]), .S0 (\genblk2.pcpi_div_n_2109
       ), .Y (n_11693));
  MXI2XL g189419(.A (\genblk2.pcpi_div_dividend [6]), .B
       (\genblk2.pcpi_div_quotient [6]), .S0 (\genblk2.pcpi_div_n_2109
       ), .Y (n_11694));
  MXI2XL g189420(.A (\genblk2.pcpi_div_dividend [8]), .B
       (\genblk2.pcpi_div_quotient [8]), .S0 (\genblk2.pcpi_div_n_2109
       ), .Y (n_11695));
  MXI2XL g189421(.A (\genblk2.pcpi_div_dividend [16]), .B
       (\genblk2.pcpi_div_quotient [16]), .S0 (\genblk2.pcpi_div_n_2109
       ), .Y (n_11696));
  MXI2XL g189422(.A (\genblk2.pcpi_div_dividend [18]), .B
       (\genblk2.pcpi_div_quotient [18]), .S0 (\genblk2.pcpi_div_n_2109
       ), .Y (n_11697));
  MXI2XL g189423(.A (\genblk2.pcpi_div_dividend [28]), .B
       (\genblk2.pcpi_div_quotient [28]), .S0 (\genblk2.pcpi_div_n_2109
       ), .Y (n_11698));
  MXI2XL g189424(.A (\genblk2.pcpi_div_dividend [22]), .B
       (\genblk2.pcpi_div_quotient [22]), .S0 (\genblk2.pcpi_div_n_2109
       ), .Y (n_11699));
  MXI2XL g189425(.A (\genblk2.pcpi_div_dividend [2]), .B
       (\genblk2.pcpi_div_quotient [2]), .S0 (\genblk2.pcpi_div_n_2109
       ), .Y (n_11700));
  MXI2XL g189426(.A (\genblk2.pcpi_div_dividend [4]), .B
       (\genblk2.pcpi_div_quotient [4]), .S0 (\genblk2.pcpi_div_n_2109
       ), .Y (n_11701));
  MXI2XL g189427(.A (\genblk2.pcpi_div_dividend [26]), .B
       (\genblk2.pcpi_div_quotient [26]), .S0 (\genblk2.pcpi_div_n_2109
       ), .Y (n_11702));
  MXI2XL g189428(.A (\genblk2.pcpi_div_dividend [20]), .B
       (\genblk2.pcpi_div_quotient [20]), .S0 (\genblk2.pcpi_div_n_2109
       ), .Y (n_11703));
  MXI2XL g189429(.A (\genblk2.pcpi_div_dividend [12]), .B
       (\genblk2.pcpi_div_quotient [12]), .S0 (\genblk2.pcpi_div_n_2109
       ), .Y (n_11704));
  MXI2XL g189430(.A (\genblk2.pcpi_div_dividend [24]), .B
       (\genblk2.pcpi_div_quotient [24]), .S0 (\genblk2.pcpi_div_n_2109
       ), .Y (n_11705));
  MXI2XL g189431(.A (\reg_op1[20]_9657 ), .B
       (\genblk2.pcpi_div_divisor [20]), .S0 (\genblk2.pcpi_div_n_4742
       ), .Y (n_11706));
  MXI2XL g189432(.A (\reg_op1[13]_9650 ), .B
       (\genblk2.pcpi_div_divisor [13]), .S0 (\genblk2.pcpi_div_n_4742
       ), .Y (n_11707));
  MXI2XL g189433(.A (\reg_op1[9]_9646 ), .B
       (\genblk2.pcpi_div_divisor [9]), .S0 (\genblk2.pcpi_div_n_4742
       ), .Y (n_11708));
  MXI2XL g189434(.A (\reg_op1[1]_9638 ), .B
       (\genblk2.pcpi_div_divisor [1]), .S0 (\genblk2.pcpi_div_n_4742
       ), .Y (n_11709));
  MXI2XL g189435(.A (\reg_op1[7]_9644 ), .B
       (\genblk2.pcpi_div_divisor [7]), .S0 (\genblk2.pcpi_div_n_4742
       ), .Y (n_11710));
  MXI2XL g189436(.A (\reg_op1[14]_9651 ), .B
       (\genblk2.pcpi_div_divisor [14]), .S0 (\genblk2.pcpi_div_n_4742
       ), .Y (n_11711));
  MXI2XL g189437(.A (\reg_op1[15]_9652 ), .B
       (\genblk2.pcpi_div_divisor [15]), .S0 (\genblk2.pcpi_div_n_4742
       ), .Y (n_11712));
  MXI2XL g189438(.A (\reg_op1[2]_9639 ), .B
       (\genblk2.pcpi_div_divisor [2]), .S0 (\genblk2.pcpi_div_n_4742
       ), .Y (n_11713));
  MXI2XL g189439(.A (\reg_op1[24]_9661 ), .B
       (\genblk2.pcpi_div_divisor [24]), .S0 (\genblk2.pcpi_div_n_4742
       ), .Y (n_11714));
  MXI2XL g189440(.A (\reg_op1[16]_9653 ), .B
       (\genblk2.pcpi_div_divisor [16]), .S0 (\genblk2.pcpi_div_n_4742
       ), .Y (n_11715));
  MXI2XL g189441(.A (\reg_op1[5]_9642 ), .B
       (\genblk2.pcpi_div_divisor [5]), .S0 (\genblk2.pcpi_div_n_4742
       ), .Y (n_11716));
  MXI2XL g189442(.A (\reg_op1[3]_9640 ), .B
       (\genblk2.pcpi_div_divisor [3]), .S0 (\genblk2.pcpi_div_n_4742
       ), .Y (n_11717));
  MXI2XL g189443(.A (\reg_op1[10]_9647 ), .B
       (\genblk2.pcpi_div_divisor [10]), .S0 (\genblk2.pcpi_div_n_4742
       ), .Y (n_11718));
  MXI2XL g189444(.A (\reg_op1[30]_9667 ), .B
       (\genblk2.pcpi_div_divisor [30]), .S0 (\genblk2.pcpi_div_n_4742
       ), .Y (n_11719));
  MXI2XL g189445(.A (\reg_op1[29]_9666 ), .B
       (\genblk2.pcpi_div_divisor [29]), .S0 (\genblk2.pcpi_div_n_4742
       ), .Y (n_11720));
  MXI2XL g189446(.A (\reg_op1[21]_9658 ), .B
       (\genblk2.pcpi_div_divisor [21]), .S0 (\genblk2.pcpi_div_n_4742
       ), .Y (n_11721));
  MXI2XL g189447(.A (\reg_op1[26]_9663 ), .B
       (\genblk2.pcpi_div_divisor [26]), .S0 (\genblk2.pcpi_div_n_4742
       ), .Y (n_11722));
  MXI2XL g189448(.A (\reg_op1[18]_9655 ), .B
       (\genblk2.pcpi_div_divisor [18]), .S0 (\genblk2.pcpi_div_n_4742
       ), .Y (n_11723));
  MXI2XL g189449(.A (\reg_op1[4]_9641 ), .B
       (\genblk2.pcpi_div_divisor [4]), .S0 (\genblk2.pcpi_div_n_4742
       ), .Y (n_11724));
  MXI2XL g189450(.A (\reg_op1[23]_9660 ), .B
       (\genblk2.pcpi_div_divisor [23]), .S0 (\genblk2.pcpi_div_n_4742
       ), .Y (n_11725));
  MXI2XL g189451(.A (\reg_op1[22]_9659 ), .B
       (\genblk2.pcpi_div_divisor [22]), .S0 (\genblk2.pcpi_div_n_4742
       ), .Y (n_11726));
  MXI2XL g189452(.A (\reg_op1[25]_9662 ), .B
       (\genblk2.pcpi_div_divisor [25]), .S0 (\genblk2.pcpi_div_n_4742
       ), .Y (n_11727));
  MXI2XL g189453(.A (\reg_op1[11]_9648 ), .B
       (\genblk2.pcpi_div_divisor [11]), .S0 (\genblk2.pcpi_div_n_4742
       ), .Y (n_11728));
  MXI2XL g189454(.A (\reg_op1[28]_9665 ), .B
       (\genblk2.pcpi_div_divisor [28]), .S0 (\genblk2.pcpi_div_n_4742
       ), .Y (n_11729));
  MXI2XL g189455(.A (\reg_op1[6]_9643 ), .B
       (\genblk2.pcpi_div_divisor [6]), .S0 (\genblk2.pcpi_div_n_4742
       ), .Y (n_11730));
  MXI2XL g189456(.A (\reg_op1[19]_9656 ), .B
       (\genblk2.pcpi_div_divisor [19]), .S0 (\genblk2.pcpi_div_n_4742
       ), .Y (n_11731));
  MXI2XL g189457(.A (\reg_op1[12]_9649 ), .B
       (\genblk2.pcpi_div_divisor [12]), .S0 (\genblk2.pcpi_div_n_4742
       ), .Y (n_11732));
  MXI2XL g189458(.A (\reg_op1[27]_9664 ), .B
       (\genblk2.pcpi_div_divisor [27]), .S0 (\genblk2.pcpi_div_n_4742
       ), .Y (n_11733));
  MXI2XL g189459(.A (\reg_op1[8]_9645 ), .B
       (\genblk2.pcpi_div_divisor [8]), .S0 (\genblk2.pcpi_div_n_4742
       ), .Y (n_11734));
  MXI2XL g189460(.A (\reg_op1[17]_9654 ), .B
       (\genblk2.pcpi_div_divisor [17]), .S0 (\genblk2.pcpi_div_n_4742
       ), .Y (n_11735));
  NOR4BX1 g189461(.AN (n_6088), .B (n_6661), .C (n_6667), .D (n_6663),
       .Y (n_11736));
  NOR4BX1 g189462(.AN (n_6090), .B (n_6671), .C (n_6665), .D (n_6666),
       .Y (n_11737));
  NOR4BBX1 g189463(.AN (n_6092), .BN (n_6091), .C (n_6668), .D
       (n_4707), .Y (n_11738));
  NAND2BX1 g189464(.AN (\reg_op1[12]_9649 ), .B (\reg_op2[12]_9681 ),
       .Y (n_11739));
  NAND2BX1 g189465(.AN (\reg_op1[13]_9650 ), .B (\reg_op2[13]_9682 ),
       .Y (n_11740));
  NAND2BX1 g189466(.AN (n_503), .B (n_440), .Y (n_11741));
  NOR2BX1 g189467(.AN (n_442), .B (latched_stalu), .Y (n_11742));
  NOR2BX1 g189468(.AN (n_425), .B (n_548), .Y (n_11743));
  NOR2BX1 g189469(.AN (n_424), .B (n_548), .Y (n_11744));
  NAND2BX1 g189470(.AN (n_338), .B (n_1335), .Y (n_11745));
  NOR2BX1 g189471(.AN (n_333), .B (n_548), .Y (n_11746));
  NOR2BX1 g189472(.AN (n_318), .B (n_1331), .Y (n_11747));
  NOR2BX1 g189473(.AN (n_291), .B (n_548), .Y (n_11748));
  NOR2BX1 g189474(.AN (n_14409_BAR), .B (n_1954), .Y (n_11749));
  NAND2BX1 g189475(.AN (\genblk1.pcpi_mul_rs2 [2]), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .Y (n_11750));
  NAND2BX1 g189476(.AN (\genblk1.pcpi_mul_rs2 [16]), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .Y (n_11751));
  NAND2BX1 g189477(.AN (\genblk1.pcpi_mul_rs2 [6]), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .Y (n_11752));
  NAND2BX1 g189478(.AN (\genblk1.pcpi_mul_rs2 [18]), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .Y (n_11753));
  NAND2BX1 g189479(.AN (\genblk1.pcpi_mul_rs2 [4]), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .Y (n_11754));
  NAND2BX1 g189480(.AN (\genblk1.pcpi_mul_rs2 [28]), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .Y (n_11755));
  NAND2BX1 g189481(.AN (\genblk1.pcpi_mul_rs2 [12]), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .Y (n_11756));
  NAND2BX1 g189482(.AN (\genblk1.pcpi_mul_rs2 [30]), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .Y (n_11757));
  NAND2BX1 g189483(.AN (\genblk1.pcpi_mul_rs2 [14]), .B
       (\genblk1.pcpi_mul_mul_2366_47_n_101 ), .Y (n_11758));
  AO22X1 g189484(.A0 (\reg_op2[24]_9693 ), .A1 (n_608), .B0
       (\reg_op2[8]_9677 ), .B1 (n_5980), .Y (n_11759));
  AO22X1 g189485(.A0 (\reg_op2[28]_9697 ), .A1 (n_608), .B0
       (\reg_op2[12]_9681 ), .B1 (n_5980), .Y (n_11760));
  AO22X1 g189486(.A0 (\reg_op2[30]_9699 ), .A1 (n_608), .B0
       (\reg_op2[14]_9683 ), .B1 (n_5980), .Y (n_11761));
  AO22X1 g189487(.A0 (\reg_op2[27]_9696 ), .A1 (n_608), .B0
       (\reg_op2[11]_9680 ), .B1 (n_5980), .Y (n_11762));
  AO22X1 g189488(.A0 (\reg_op2[31]_9700 ), .A1 (n_608), .B0
       (\reg_op2[15]_9684 ), .B1 (n_5980), .Y (n_11763));
  AO22X1 g189489(.A0 (\reg_op2[26]_9695 ), .A1 (n_608), .B0
       (\reg_op2[10]_9679 ), .B1 (n_5980), .Y (n_11764));
  AO22X1 g189490(.A0 (\reg_op2[29]_9698 ), .A1 (n_608), .B0
       (\reg_op2[13]_9682 ), .B1 (n_5980), .Y (n_11765));
  AO22X1 g189491(.A0 (\reg_op2[25]_9694 ), .A1 (n_608), .B0
       (\reg_op2[9]_9678 ), .B1 (n_5980), .Y (n_11766));
  AO22X1 g189492(.A0 (\genblk2.pcpi_div_quotient_msk [31]), .A1
       (n_444), .B0 (\genblk2.pcpi_div_quotient [31]), .B1 (n_954), .Y
       (n_11767));
  AO22X1 g189493(.A0 (\genblk2.pcpi_div_quotient_msk [0]), .A1 (n_444),
       .B0 (\genblk2.pcpi_div_quotient [0]), .B1 (n_954), .Y (n_11768));
  AO22X1 g189494(.A0 (\genblk2.pcpi_div_quotient_msk [1]), .A1 (n_444),
       .B0 (\genblk2.pcpi_div_quotient [1]), .B1 (n_954), .Y (n_11769));
  AO22X1 g189495(.A0 (\genblk2.pcpi_div_quotient_msk [2]), .A1 (n_444),
       .B0 (\genblk2.pcpi_div_quotient [2]), .B1 (n_954), .Y (n_11770));
  AO22X1 g189496(.A0 (\genblk2.pcpi_div_quotient_msk [3]), .A1 (n_444),
       .B0 (\genblk2.pcpi_div_quotient [3]), .B1 (n_954), .Y (n_11771));
  AO22X1 g189497(.A0 (\genblk2.pcpi_div_quotient_msk [4]), .A1 (n_444),
       .B0 (\genblk2.pcpi_div_quotient [4]), .B1 (n_954), .Y (n_11772));
  AO22X1 g189498(.A0 (\genblk2.pcpi_div_quotient_msk [5]), .A1 (n_444),
       .B0 (\genblk2.pcpi_div_quotient [5]), .B1 (n_954), .Y (n_11773));
  AO22X1 g189499(.A0 (\genblk2.pcpi_div_quotient_msk [7]), .A1 (n_444),
       .B0 (\genblk2.pcpi_div_quotient [7]), .B1 (n_954), .Y (n_11774));
  AO22X1 g189500(.A0 (\genblk2.pcpi_div_quotient_msk [6]), .A1 (n_444),
       .B0 (\genblk2.pcpi_div_quotient [6]), .B1 (n_954), .Y (n_11775));
  AO22X1 g189501(.A0 (\genblk2.pcpi_div_quotient_msk [8]), .A1 (n_444),
       .B0 (\genblk2.pcpi_div_quotient [8]), .B1 (n_954), .Y (n_11776));
  AO22X1 g189502(.A0 (\genblk2.pcpi_div_quotient_msk [9]), .A1 (n_444),
       .B0 (\genblk2.pcpi_div_quotient [9]), .B1 (n_954), .Y (n_11777));
  AO22X1 g189503(.A0 (\genblk2.pcpi_div_quotient_msk [10]), .A1
       (n_444), .B0 (\genblk2.pcpi_div_quotient [10]), .B1 (n_954), .Y
       (n_11778));
  AO22X1 g189504(.A0 (\genblk2.pcpi_div_quotient_msk [11]), .A1
       (n_444), .B0 (\genblk2.pcpi_div_quotient [11]), .B1 (n_954), .Y
       (n_11779));
  AO22X1 g189505(.A0 (\genblk2.pcpi_div_quotient_msk [12]), .A1
       (n_444), .B0 (\genblk2.pcpi_div_quotient [12]), .B1 (n_954), .Y
       (n_11780));
  AO22X1 g189506(.A0 (\genblk2.pcpi_div_quotient_msk [13]), .A1
       (n_444), .B0 (\genblk2.pcpi_div_quotient [13]), .B1 (n_954), .Y
       (n_11781));
  AO22X1 g189507(.A0 (\genblk2.pcpi_div_quotient_msk [14]), .A1
       (n_444), .B0 (\genblk2.pcpi_div_quotient [14]), .B1 (n_954), .Y
       (n_11782));
  AO22X1 g189508(.A0 (\genblk2.pcpi_div_quotient_msk [15]), .A1
       (n_444), .B0 (\genblk2.pcpi_div_quotient [15]), .B1 (n_954), .Y
       (n_11783));
  AO22X1 g189509(.A0 (\genblk2.pcpi_div_quotient_msk [16]), .A1
       (n_444), .B0 (\genblk2.pcpi_div_quotient [16]), .B1 (n_954), .Y
       (n_11784));
  AO22X1 g189510(.A0 (\genblk2.pcpi_div_quotient_msk [17]), .A1
       (n_444), .B0 (\genblk2.pcpi_div_quotient [17]), .B1 (n_954), .Y
       (n_11785));
  AO22X1 g189511(.A0 (\genblk2.pcpi_div_quotient_msk [18]), .A1
       (n_444), .B0 (\genblk2.pcpi_div_quotient [18]), .B1 (n_954), .Y
       (n_11786));
  AO22X1 g189512(.A0 (\genblk2.pcpi_div_quotient_msk [19]), .A1
       (n_444), .B0 (\genblk2.pcpi_div_quotient [19]), .B1 (n_954), .Y
       (n_11787));
  AO22X1 g189513(.A0 (\genblk2.pcpi_div_quotient_msk [20]), .A1
       (n_444), .B0 (\genblk2.pcpi_div_quotient [20]), .B1 (n_954), .Y
       (n_11788));
  AO22X1 g189514(.A0 (\genblk2.pcpi_div_quotient_msk [22]), .A1
       (n_444), .B0 (\genblk2.pcpi_div_quotient [22]), .B1 (n_954), .Y
       (n_11789));
  AO22X1 g189515(.A0 (\genblk2.pcpi_div_quotient_msk [23]), .A1
       (n_444), .B0 (\genblk2.pcpi_div_quotient [23]), .B1 (n_954), .Y
       (n_11790));
  AO22X1 g189516(.A0 (\genblk2.pcpi_div_quotient_msk [21]), .A1
       (n_444), .B0 (\genblk2.pcpi_div_quotient [21]), .B1 (n_954), .Y
       (n_11791));
  AO22X1 g189517(.A0 (\genblk2.pcpi_div_quotient_msk [24]), .A1
       (n_444), .B0 (\genblk2.pcpi_div_quotient [24]), .B1 (n_954), .Y
       (n_11792));
  AO22X1 g189518(.A0 (\genblk2.pcpi_div_quotient_msk [25]), .A1
       (n_444), .B0 (\genblk2.pcpi_div_quotient [25]), .B1 (n_954), .Y
       (n_11793));
  AO22X1 g189519(.A0 (\genblk2.pcpi_div_quotient_msk [26]), .A1
       (n_444), .B0 (\genblk2.pcpi_div_quotient [26]), .B1 (n_954), .Y
       (n_11794));
  AO22X1 g189520(.A0 (\genblk2.pcpi_div_quotient_msk [27]), .A1
       (n_444), .B0 (\genblk2.pcpi_div_quotient [27]), .B1 (n_954), .Y
       (n_11795));
  AO22X1 g189521(.A0 (\genblk2.pcpi_div_quotient_msk [28]), .A1
       (n_444), .B0 (\genblk2.pcpi_div_quotient [28]), .B1 (n_954), .Y
       (n_11796));
  AO22X1 g189522(.A0 (\genblk2.pcpi_div_quotient_msk [29]), .A1
       (n_444), .B0 (\genblk2.pcpi_div_quotient [29]), .B1 (n_954), .Y
       (n_11797));
  AO22X1 g189523(.A0 (\genblk2.pcpi_div_quotient_msk [30]), .A1
       (n_444), .B0 (\genblk2.pcpi_div_quotient [30]), .B1 (n_954), .Y
       (n_11798));
  AO22X1 g189524(.A0 (n_446), .A1 (n_437), .B0 (mem_rdata_q[3]), .B1
       (n_445), .Y (n_11799));
  AO22X1 g189525(.A0 (\cpuregs[25] [0]), .A1 (n_1594), .B0
       (\cpuregs[26] [0]), .B1 (n_1613), .Y (n_11800));
  AO22X1 g189526(.A0 (reg_pc[16]), .A1 (n_427), .B0 (current_pc[16]),
       .B1 (n_658), .Y (n_11801));
  AO22X1 g189527(.A0 (reg_pc[9]), .A1 (n_427), .B0 (current_pc[9]), .B1
       (n_658), .Y (n_11802));
  AO22X1 g189528(.A0 (reg_pc[8]), .A1 (n_427), .B0 (current_pc[8]), .B1
       (n_658), .Y (n_11803));
  AO22X1 g189529(.A0 (reg_pc[25]), .A1 (n_427), .B0 (current_pc[25]),
       .B1 (n_658), .Y (n_11804));
  AO22X1 g189530(.A0 (reg_pc[17]), .A1 (n_427), .B0 (current_pc[17]),
       .B1 (n_658), .Y (n_11805));
  AO22X1 g189531(.A0 (reg_pc[24]), .A1 (n_427), .B0 (current_pc[24]),
       .B1 (n_658), .Y (n_11806));
  AO22X1 g189532(.A0 (reg_pc[15]), .A1 (n_427), .B0 (current_pc[15]),
       .B1 (n_658), .Y (n_11807));
  AO22X1 g189533(.A0 (reg_pc[28]), .A1 (n_427), .B0 (current_pc[28]),
       .B1 (n_658), .Y (n_11808));
  AO22X1 g189534(.A0 (reg_pc[19]), .A1 (n_427), .B0 (current_pc[19]),
       .B1 (n_658), .Y (n_11809));
  AO22X1 g189535(.A0 (reg_pc[20]), .A1 (n_427), .B0 (current_pc[20]),
       .B1 (n_658), .Y (n_11810));
  AO22X1 g189536(.A0 (reg_pc[29]), .A1 (n_427), .B0 (current_pc[29]),
       .B1 (n_658), .Y (n_11811));
  AO22X1 g189537(.A0 (reg_pc[12]), .A1 (n_427), .B0 (current_pc[12]),
       .B1 (n_658), .Y (n_11812));
  AO22X1 g189538(.A0 (reg_pc[21]), .A1 (n_427), .B0 (current_pc[21]),
       .B1 (n_658), .Y (n_11813));
  AO22X1 g189539(.A0 (reg_pc[14]), .A1 (n_427), .B0 (current_pc[14]),
       .B1 (n_658), .Y (n_11814));
  AO22X1 g189540(.A0 (reg_pc[31]), .A1 (n_427), .B0 (current_pc[31]),
       .B1 (n_658), .Y (n_11815));
  AO22X1 g189541(.A0 (reg_pc[23]), .A1 (n_427), .B0 (current_pc[23]),
       .B1 (n_658), .Y (n_11816));
  AO22X1 g189542(.A0 (reg_pc[13]), .A1 (n_427), .B0 (current_pc[13]),
       .B1 (n_658), .Y (n_11817));
  AO22X1 g189543(.A0 (reg_pc[27]), .A1 (n_427), .B0 (current_pc[27]),
       .B1 (n_658), .Y (n_11818));
  AO22X1 g189544(.A0 (reg_pc[18]), .A1 (n_427), .B0 (current_pc[18]),
       .B1 (n_658), .Y (n_11819));
  AO22X1 g189545(.A0 (reg_pc[10]), .A1 (n_427), .B0 (current_pc[10]),
       .B1 (n_658), .Y (n_11820));
  AO22X1 g189546(.A0 (reg_pc[2]), .A1 (n_427), .B0 (current_pc[2]), .B1
       (n_658), .Y (n_11821));
  AO22X1 g189547(.A0 (reg_pc[5]), .A1 (n_427), .B0 (current_pc[5]), .B1
       (n_658), .Y (n_11822));
  AO22X1 g189548(.A0 (reg_pc[4]), .A1 (n_427), .B0 (current_pc[4]), .B1
       (n_658), .Y (n_11823));
  AO22X1 g189549(.A0 (reg_pc[6]), .A1 (n_427), .B0 (current_pc[6]), .B1
       (n_658), .Y (n_11824));
  AO22X1 g189550(.A0 (reg_pc[3]), .A1 (n_427), .B0 (current_pc[3]), .B1
       (n_658), .Y (n_11825));
  AO22X1 g189551(.A0 (reg_pc[1]), .A1 (n_427), .B0 (current_pc[1]), .B1
       (n_658), .Y (n_11826));
  AO22X1 g189552(.A0 (reg_pc[11]), .A1 (n_427), .B0 (current_pc[11]),
       .B1 (n_658), .Y (n_11827));
  AO22X1 g189553(.A0 (reg_pc[26]), .A1 (n_427), .B0 (current_pc[26]),
       .B1 (n_658), .Y (n_11828));
  AO22X1 g189554(.A0 (reg_pc[30]), .A1 (n_427), .B0 (current_pc[30]),
       .B1 (n_658), .Y (n_11829));
  AO22X1 g189555(.A0 (reg_pc[22]), .A1 (n_427), .B0 (current_pc[22]),
       .B1 (n_658), .Y (n_11830));
  AO22X1 g189556(.A0 (reg_pc[7]), .A1 (n_427), .B0 (current_pc[7]), .B1
       (n_658), .Y (n_11831));
  AO21X1 g189558(.A0 (n_6828), .A1 (n_313), .B0 (n_61806_BAR), .Y
       (n_11833));
  AO21X1 g189559(.A0 (n_6827), .A1 (n_313), .B0 (n_61804_BAR), .Y
       (n_11834));
  AO21X1 g189561(.A0 (n_6824), .A1 (n_313), .B0 (n_61798_BAR), .Y
       (n_11836));
  AO21X1 g189563(.A0 (n_6821), .A1 (n_313), .B0 (n_61792_BAR), .Y
       (n_11838));
  AO21X1 g189565(.A0 (n_6817), .A1 (n_313), .B0 (n_61784_BAR), .Y
       (n_11840));
  AO21X1 g189567(.A0 (n_6803), .A1 (n_313), .B0 (n_61756_BAR), .Y
       (n_11842));
  AO21X1 g189568(.A0 (n_5984), .A1 (\reg_op2[10]_9679 ), .B0 (n_6103),
       .Y (n_11843));
  AO21X1 g189569(.A0 (n_5984), .A1 (\reg_op2[14]_9683 ), .B0 (n_6141),
       .Y (n_11844));
  AO21X1 g189570(.A0 (n_6806), .A1 (n_313), .B0 (n_61762_BAR), .Y
       (n_11845));
  AO21X1 g189571(.A0 (n_6805), .A1 (n_313), .B0 (n_61760_BAR), .Y
       (n_11846));
  AO21X1 g189572(.A0 (n_6804), .A1 (n_313), .B0 (n_61758_BAR), .Y
       (n_11847));
  AO21X1 g189573(.A0 (n_5984), .A1 (\reg_op2[15]_9684 ), .B0 (n_6105),
       .Y (n_11848));
  AO21X1 g189574(.A0 (n_5984), .A1 (\reg_op2[13]_9682 ), .B0 (n_6098),
       .Y (n_11849));
  AO21X1 g189575(.A0 (n_5984), .A1 (\reg_op2[12]_9681 ), .B0 (n_6104),
       .Y (n_11850));
  AO21X1 g189576(.A0 (n_5984), .A1 (\reg_op2[11]_9680 ), .B0 (n_6101),
       .Y (n_11851));
  AO21X1 g189577(.A0 (n_5984), .A1 (\reg_op2[9]_9678 ), .B0 (n_6097),
       .Y (n_11852));
  AO21X1 g189578(.A0 (n_5984), .A1 (\reg_op2[8]_9677 ), .B0 (n_6134),
       .Y (n_11853));
  MXI2XL g189579(.A (n_5788), .B (n_11854), .S0 (n_313), .Y (n_11855));
  OAI21X1 g189580(.A0 (n_6859), .A1 (inc_add_382_74_n_222), .B0
       (inc_add_382_74_n_217), .Y (n_11854));
  MXI2XL g189581(.A (n_713), .B (n_11856), .S0 (n_313), .Y (n_11857));
  OAI21X1 g189582(.A0 (n_6855), .A1 (inc_add_382_74_n_242), .B0
       (inc_add_382_74_n_237), .Y (n_11856));
  MXI2XL g189583(.A (n_637), .B (n_11858), .S0 (n_313), .Y (n_11859));
  OAI21X1 g189584(.A0 (n_6852), .A1 (inc_add_382_74_n_257), .B0
       (inc_add_382_74_n_252), .Y (n_11858));
  MXI2XL g189585(.A (n_715), .B (n_11860), .S0 (n_313), .Y (n_11861));
  OAI21X1 g189586(.A0 (n_6848), .A1 (inc_add_382_74_n_277), .B0
       (inc_add_382_74_n_272), .Y (n_11860));
  MXI2XL g189587(.A (n_718), .B (n_11862), .S0 (n_313), .Y (n_11863));
  OAI21X1 g189588(.A0 (n_6861), .A1 (inc_add_382_74_n_212), .B0
       (inc_add_382_74_n_207), .Y (n_11862));
  AND2X1 g190057(.A (n_6514), .B (n_538), .Y (n_13034));
endmodule

module picorv32_chip(clk, resetn, trap, mem_valid, mem_instr, mem_ready,
     mem_addr, mem_wdata, mem_wstrb, mem_rdata, mem_la_read,
     mem_la_write, mem_la_addr, mem_la_wdata, mem_la_wstrb, pcpi_valid,
     pcpi_insn, pcpi_rs1, pcpi_rs2, pcpi_wr, pcpi_rd, pcpi_wait,
     pcpi_ready, irq, eoi, trace_valid, trace_data);

     input clk, resetn, mem_ready, pcpi_wr, pcpi_wait, pcpi_ready;
     input [31:0] mem_rdata, pcpi_rd, irq;
     output trap, mem_valid, mem_instr, mem_la_read, mem_la_write,
          pcpi_valid, trace_valid;
     output [31:0] mem_addr, mem_wdata, mem_la_addr, mem_la_wdata,
          pcpi_insn, pcpi_rs1, pcpi_rs2, eoi;
     output [3:0] mem_wstrb, mem_la_wstrb;
     output [35:0] trace_data;
     wire clk_w, resetn_w, mem_ready_w, pcpi_wr_w, pcpi_wait_w, pcpi_ready_w;
     wire [31:0] mem_rdata_w, pcpi_rd_w, irq_w;
     wire trap_w, mem_valid_w, mem_instr_w, mem_la_read_w, mem_la_write_w,
          pcpi_valid_w, trace_valid_w;
     wire [31:0] mem_addr_w, mem_wdata_w, mem_la_addr_w, mem_la_wdata_w,
          pcpi_insn_w, pcpi_rs1_w, pcpi_rs2_w, eoi_w;
     wire [3:0] mem_wstrb_w, mem_la_wstrb_w;
     wire [35:0] trace_data_w;

     picorv32 example(clk_w, resetn_w, trap_w, mem_valid_w, mem_instr_w, mem_ready_w,
     mem_addr_w, mem_wdata_w, mem_wstrb_w, mem_rdata_w, mem_la_read_w,
     mem_la_write_w, mem_la_addr_w, mem_la_wdata_w, mem_la_wstrb_w, pcpi_valid_w,
     pcpi_insn_w, pcpi_rs1_w, pcpi_rs2_w, pcpi_wr_w, pcpi_rd_w, pcpi_wait_w,
     pcpi_ready_w, irq_w, eoi_w, trace_valid_w, trace_data_w);
  
 picorv32_pads iopads(clk, resetn, trap, mem_valid, mem_instr, mem_ready,
     mem_addr, mem_wdata, mem_wstrb, mem_rdata, mem_la_read,
     mem_la_write, mem_la_addr, mem_la_wdata, mem_la_wstrb, pcpi_valid,
     pcpi_insn, pcpi_rs1, pcpi_rs2, pcpi_wr, pcpi_rd, pcpi_wait,
     pcpi_ready, irq, eoi, trace_valid, trace_data, 
     clk_w, resetn_w, trap_w, mem_valid_w, mem_instr_w, mem_ready_w,
     mem_addr_w, mem_wdata_w, mem_wstrb_w, mem_rdata_w, mem_la_read_w,
     mem_la_write_w, mem_la_addr_w, mem_la_wdata_w, mem_la_wstrb_w, pcpi_valid_w,
     pcpi_insn_w, pcpi_rs1_w, pcpi_rs2_w, pcpi_wr_w, pcpi_rd_w, pcpi_wait_w,
     pcpi_ready_w, irq_w, eoi_w, trace_valid_w, trace_data_w, VSS, VDD);
endmodule


